//------------------------------------------------------------------------------
// The confidential and proprietary information contained in this file may
// only be used by a person authorised under and to the extent permitted
// by a subsisting licensing agreement from ARM Limited.
//
//            (C) COPYRIGHT 2010 ARM Limited.
//                ALL RIGHTS RESERVED
//
// This entire notice must be reproduced on all copies of this file
// and copies of this file may only be made by a person if such person is
// permitted to do so under the terms of a subsisting license agreement
// from ARM Limited.
//
//      SVN Information
//
//      Checked In          : 2010-08-03 21:05:56 +0100 (Tue, 03 Aug 2010)
//
//      Revision            : 144987
//
//      Release Information : AT510-MN-80001-r0p0-00rel0
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Cortex-M0 DesignStart processor logic level
//------------------------------------------------------------------------------

module cortexm0ds_logic
(hclk, hreset_n, haddr_o, hburst_o, hmastlock_o, hprot_o,
hsize_o, htrans_o, hwdata_o, hwrite_o, hrdata_i, hready_i, hresp_i,
nmi_i, irq_i, txev_o, rxev_i, lockup_o, sys_reset_req_o, sleeping_o,
vis_r0_o, vis_r1_o, vis_r2_o, vis_r3_o, vis_r4_o, vis_r5_o, vis_r6_o,
vis_r7_o, vis_r8_o, vis_r9_o, vis_r10_o, vis_r11_o, vis_r12_o, vis_r14_o
, vis_msp_o, vis_psp_o, vis_pc_o, vis_apsr_o, vis_tbit_o, vis_ipsr_o,
vis_control_o, vis_primask_o);

output [31:0] haddr_o;
output [2:0] hburst_o;
output [3:0] hprot_o;
output [2:0] hsize_o;
output [1:0] htrans_o;
output [31:0] hwdata_o;
input [31:0] hrdata_i;
input [15:0] irq_i;
output [31:0] vis_r0_o;
output [31:0] vis_r1_o;
output [31:0] vis_r2_o;
output [31:0] vis_r3_o;
output [31:0] vis_r4_o;
output [31:0] vis_r5_o;
output [31:0] vis_r6_o;
output [31:0] vis_r7_o;
output [31:0] vis_r8_o;
output [31:0] vis_r9_o;
output [31:0] vis_r10_o;
output [31:0] vis_r11_o;
output [31:0] vis_r12_o;
output [31:0] vis_r14_o;
output [29:0] vis_msp_o;
output [29:0] vis_psp_o;
output [30:0] vis_pc_o;
output [3:0] vis_apsr_o;
output [5:0] vis_ipsr_o;
input hclk;
input hreset_n;
input hready_i;
input hresp_i;
input nmi_i;
input rxev_i;
output hmastlock_o;
output hwrite_o;
output txev_o;
output lockup_o;
output sys_reset_req_o;
output sleeping_o;
output vis_tbit_o;
output vis_control_o;
output vis_primask_o;

wire Mf8vx4, Eg8vx4, Ih8vx4, Ki8vx4, Mj8vx4, Mk8vx4, Ul8vx4, Cn8vx4, Ho8vx4, Pp8vx4;
wire Xq8vx4, Fs8vx4, Nt8vx4, Vu8vx4, Dw8vx4, Hx8vx4, Oy8vx4, Uz8vx4, B19vx4, I29vx4;
wire P39vx4, W49vx4, D69vx4, K79vx4, R89vx4, Y99vx4, Fb9vx4, Mc9vx4, Ud9vx4, Cf9vx4;
wire Kg9vx4, Sh9vx4, Aj9vx4, Ik9vx4, Ml9vx4, Qm9vx4, Un9vx4, Yo9vx4, Cq9vx4, Gr9vx4;
wire Ks9vx4, Ot9vx4, Su9vx4, Wv9vx4, Bx9vx4, Gy9vx4, Jz9vx4, M0avx4, P1avx4, S2avx4;
wire V3avx4, Y4avx4, B6avx4, E7avx4, H8avx4, K9avx4, Naavx4, Qbavx4, Tcavx4, Wdavx4;
wire Zeavx4, Cgavx4, Fhavx4, Iiavx4, Ljavx4, Okavx4, Rlavx4, Umavx4, Xnavx4, Apavx4;
wire Dqavx4, Gravx4, Jsavx4, Ltavx4, Nuavx4, Pvavx4, Rwavx4, Txavx4, Vyavx4, Xzavx4;
wire E1bvx4, O2bvx4, Y3bvx4, I5bvx4, T6bvx4, E8bvx4, P9bvx4, Abbvx4, Lcbvx4, Wdbvx4;
wire Hfbvx4, Sgbvx4, Dibvx4, Ojbvx4, Zkbvx4, Kmbvx4, Vnbvx4, Gpbvx4, Qqbvx4, Asbvx4;
wire Ktbvx4, Uubvx4, Ewbvx4, Oxbvx4, Yybvx4, I0cvx4, S1cvx4, C3cvx4, N4cvx4, Y5cvx4;
wire J7cvx4, U8cvx4, Facvx4, Qbcvx4, Bdcvx4, Mecvx4, Xfcvx4, Ihcvx4, Ticvx4, Ekcvx4;
wire Plcvx4, Ancvx4, Locvx4, Wpcvx4, Hrcvx4, Sscvx4, Ducvx4, Ovcvx4, Zwcvx4, Kycvx4;
wire Uzcvx4, E1dvx4, O2dvx4, Y3dvx4, I5dvx4, S6dvx4, C8dvx4, M9dvx4, Wadvx4, Gcdvx4;
wire Rddvx4, Cfdvx4, Ngdvx4, Yhdvx4, Jjdvx4, Ukdvx4, Fmdvx4, Qndvx4, Bpdvx4, Mqdvx4;
wire Xrdvx4, Itdvx4, Tudvx4, Ewdvx4, Pxdvx4, Azdvx4, L0evx4, W1evx4, H3evx4, S4evx4;
wire D6evx4, O7evx4, V8evx4, Faevx4, Rbevx4, Ddevx4, Peevx4, Bgevx4, Nhevx4, Zievx4;
wire Lkevx4, Xlevx4, Hnevx4, Roevx4, Bqevx4, Lrevx4, Vsevx4, Fuevx4, Pvevx4, Zwevx4;
wire Jyevx4, Tzevx4, D1fvx4, O2fvx4, Z3fvx4, K5fvx4, V6fvx4, G8fvx4, R9fvx4, Cbfvx4;
wire Mcfvx4, Wdfvx4, Gffvx4, Qgfvx4, Aifvx4, Kjfvx4, Ukfvx4, Emfvx4, Onfvx4, Yofvx4;
wire Jqfvx4, Urfvx4, Ftfvx4, Qufvx4, Bwfvx4, Mxfvx4, Xyfvx4, H0gvx4, P1gvx4, A3gvx4;
wire I4gvx4, Q5gvx4, Z6gvx4, O8gvx4, U9gvx4, Dbgvx4, Mcgvx4, Vdgvx4, Efgvx4, Nggvx4;
wire Whgvx4, Fjgvx4, Rkgvx4, Dmgvx4, Nngvx4, Vogvx4, Eqgvx4, Krgvx4, Qsgvx4, Wtgvx4;
wire Cvgvx4, Owgvx4, Aygvx4, Izgvx4, S0hvx4, F2hvx4, R3hvx4, B5hvx4, N6hvx4, Z7hvx4;
wire L9hvx4, Xahvx4, Jchvx4, Qchvx4, Xchvx4, Edhvx4, Ldhvx4, Sdhvx4, Zdhvx4, Gehvx4;
wire Nehvx4, Uehvx4, Bfhvx4, Ifhvx4, Pfhvx4, Wfhvx4, Dghvx4, Kghvx4, Rghvx4, Yghvx4;
wire Fhhvx4, Mhhvx4, Thhvx4, Aihvx4, Hihvx4, Oihvx4, Vihvx4, Cjhvx4, Jjhvx4, Qjhvx4;
wire Xjhvx4, Ekhvx4, Lkhvx4, Skhvx4, Zkhvx4, Glhvx4, Nlhvx4, Ulhvx4, Bmhvx4, Imhvx4;
wire Pmhvx4, Wmhvx4, Dnhvx4, Knhvx4, Rnhvx4, Ynhvx4, Fohvx4, Mohvx4, Tohvx4, Aphvx4;
wire Hphvx4, Ophvx4, Vphvx4, Cqhvx4, Jqhvx4, Qqhvx4, Xqhvx4, Erhvx4, Lrhvx4, Srhvx4;
wire Zrhvx4, Gshvx4, Nshvx4, Ushvx4, Bthvx4, Ithvx4, Pthvx4, Wthvx4, Duhvx4, Kuhvx4;
wire Ruhvx4, Yuhvx4, Fvhvx4, Mvhvx4, Tvhvx4, Awhvx4, Hwhvx4, Owhvx4, Vwhvx4, Cxhvx4;
wire Jxhvx4, Qxhvx4, Xxhvx4, Eyhvx4, Lyhvx4, Syhvx4, Zyhvx4, Gzhvx4, Nzhvx4, Uzhvx4;
wire B0ivx4, I0ivx4, P0ivx4, W0ivx4, D1ivx4, K1ivx4, R1ivx4, Y1ivx4, F2ivx4, M2ivx4;
wire T2ivx4, A3ivx4, H3ivx4, O3ivx4, V3ivx4, C4ivx4, J4ivx4, Q4ivx4, X4ivx4, E5ivx4;
wire L5ivx4, S5ivx4, Z5ivx4, G6ivx4, N6ivx4, U6ivx4, B7ivx4, I7ivx4, P7ivx4, W7ivx4;
wire D8ivx4, K8ivx4, R8ivx4, Y8ivx4, F9ivx4, M9ivx4, T9ivx4, Aaivx4, Haivx4, Oaivx4;
wire Vaivx4, Cbivx4, Jbivx4, Qbivx4, Xbivx4, Ecivx4, Lcivx4, Scivx4, Zcivx4, Gdivx4;
wire Ndivx4, Udivx4, Beivx4, Ieivx4, Peivx4, Weivx4, Dfivx4, Kfivx4, Rfivx4, Yfivx4;
wire Fgivx4, Mgivx4, Tgivx4, Ahivx4, Hhivx4, Ohivx4, Vhivx4, Ciivx4, Jiivx4, Qiivx4;
wire Xiivx4, Ejivx4, Ljivx4, Sjivx4, Zjivx4, Gkivx4, Nkivx4, Ukivx4, Blivx4, Ilivx4;
wire Plivx4, Wlivx4, Dmivx4, Kmivx4, Rmivx4, Ymivx4, Fnivx4, Mnivx4, Tnivx4, Aoivx4;
wire Hoivx4, Ooivx4, Voivx4, Cpivx4, Jpivx4, Qpivx4, Xpivx4, Eqivx4, Lqivx4, Sqivx4;
wire Zqivx4, Grivx4, Nrivx4, Urivx4, Bsivx4, Isivx4, Psivx4, Wsivx4, Dtivx4, Ktivx4;
wire Rtivx4, Ytivx4, Fuivx4, Muivx4, Tuivx4, Avivx4, Hvivx4, Ovivx4, Vvivx4, Cwivx4;
wire Jwivx4, Qwivx4, Xwivx4, Exivx4, Lxivx4, Sxivx4, Zxivx4, Gyivx4, Nyivx4, Uyivx4;
wire Bzivx4, Izivx4, Pzivx4, Wzivx4, D0jvx4, K0jvx4, R0jvx4, Y0jvx4, F1jvx4, M1jvx4;
wire T1jvx4, A2jvx4, H2jvx4, O2jvx4, V2jvx4, C3jvx4, J3jvx4, Q3jvx4, X3jvx4, E4jvx4;
wire L4jvx4, S4jvx4, Z4jvx4, G5jvx4, N5jvx4, U5jvx4, B6jvx4, I6jvx4, P6jvx4, W6jvx4;
wire D7jvx4, K7jvx4, R7jvx4, Y7jvx4, F8jvx4, M8jvx4, T8jvx4, A9jvx4, H9jvx4, O9jvx4;
wire V9jvx4, Cajvx4, Jajvx4, Qajvx4, Xajvx4, Ebjvx4, Lbjvx4, Sbjvx4, Zbjvx4, Gcjvx4;
wire Ncjvx4, Ucjvx4, Bdjvx4, Idjvx4, Pdjvx4, Wdjvx4, Dejvx4, Kejvx4, Rejvx4, Yejvx4;
wire Ffjvx4, Mfjvx4, Tfjvx4, Agjvx4, Hgjvx4, Ogjvx4, Vgjvx4, Chjvx4, Jhjvx4, Qhjvx4;
wire Xhjvx4, Eijvx4, Lijvx4, Sijvx4, Zijvx4, Gjjvx4, Njjvx4, Ujjvx4, Bkjvx4, Ikjvx4;
wire Pkjvx4, Wkjvx4, Dljvx4, Kljvx4, Rljvx4, Yljvx4, Fmjvx4, Mmjvx4, Tmjvx4, Anjvx4;
wire Hnjvx4, Onjvx4, Vnjvx4, Cojvx4, Jojvx4, Qojvx4, Xojvx4, Epjvx4, Lpjvx4, Spjvx4;
wire Zpjvx4, Gqjvx4, Nqjvx4, Uqjvx4, Brjvx4, Irjvx4, Prjvx4, Wrjvx4, Dsjvx4, Ksjvx4;
wire Rsjvx4, Ysjvx4, Ftjvx4, Mtjvx4, Ttjvx4, Aujvx4, Hujvx4, Oujvx4, Vujvx4, Cvjvx4;
wire Jvjvx4, Qvjvx4, Xvjvx4, Ewjvx4, Lwjvx4, Swjvx4, Zwjvx4, Gxjvx4, Nxjvx4, Uxjvx4;
wire Byjvx4, Iyjvx4, Pyjvx4, Wyjvx4, Dzjvx4, Kzjvx4, Rzjvx4, Yzjvx4, F0kvx4, M0kvx4;
wire T0kvx4, A1kvx4, H1kvx4, O1kvx4, V1kvx4, C2kvx4, J2kvx4, Q2kvx4, X2kvx4, E3kvx4;
wire L3kvx4, S3kvx4, Z3kvx4, G4kvx4, N4kvx4, U4kvx4, B5kvx4, I5kvx4, P5kvx4, W5kvx4;
wire D6kvx4, K6kvx4, R6kvx4, Y6kvx4, F7kvx4, M7kvx4, T7kvx4, A8kvx4, H8kvx4, O8kvx4;
wire V8kvx4, C9kvx4, J9kvx4, Q9kvx4, X9kvx4, Eakvx4, Lakvx4, Sakvx4, Zakvx4, Gbkvx4;
wire Nbkvx4, Ubkvx4, Bckvx4, Ickvx4, Pckvx4, Wckvx4, Ddkvx4, Kdkvx4, Rdkvx4, Ydkvx4;
wire Fekvx4, Mekvx4, Tekvx4, Afkvx4, Hfkvx4, Ofkvx4, Vfkvx4, Cgkvx4, Jgkvx4, Qgkvx4;
wire Xgkvx4, Ehkvx4, Lhkvx4, Shkvx4, Zhkvx4, Gikvx4, Nikvx4, Uikvx4, Bjkvx4, Ijkvx4;
wire Pjkvx4, Wjkvx4, Dkkvx4, Kkkvx4, Rkkvx4, Ykkvx4, Flkvx4, Mlkvx4, Tlkvx4, Amkvx4;
wire Hmkvx4, Omkvx4, Vmkvx4, Cnkvx4, Jnkvx4, Qnkvx4, Xnkvx4, Eokvx4, Lokvx4, Sokvx4;
wire Zokvx4, Gpkvx4, Npkvx4, Upkvx4, Bqkvx4, Iqkvx4, Pqkvx4, Wqkvx4, Drkvx4, Krkvx4;
wire Rrkvx4, Yrkvx4, Fskvx4, Mskvx4, Tskvx4, Atkvx4, Htkvx4, Otkvx4, Vtkvx4, Cukvx4;
wire Jukvx4, Qukvx4, Xukvx4, Evkvx4, Lvkvx4, Svkvx4, Zvkvx4, Gwkvx4, Nwkvx4, Uwkvx4;
wire Bxkvx4, Ixkvx4, Pxkvx4, Wxkvx4, Dykvx4, Kykvx4, Rykvx4, Yykvx4, Fzkvx4, Mzkvx4;
wire Tzkvx4, A0lvx4, H0lvx4, O0lvx4, V0lvx4, C1lvx4, J1lvx4, Q1lvx4, X1lvx4, E2lvx4;
wire L2lvx4, S2lvx4, Z2lvx4, G3lvx4, N3lvx4, U3lvx4, B4lvx4, I4lvx4, P4lvx4, W4lvx4;
wire D5lvx4, K5lvx4, R5lvx4, Y5lvx4, F6lvx4, M6lvx4, T6lvx4, A7lvx4, H7lvx4, O7lvx4;
wire V7lvx4, C8lvx4, J8lvx4, Q8lvx4, X8lvx4, E9lvx4, L9lvx4, S9lvx4, Z9lvx4, Galvx4;
wire Nalvx4, Ualvx4, Bblvx4, Iblvx4, Pblvx4, Wblvx4, Dclvx4, Kclvx4, Rclvx4, Yclvx4;
wire Fdlvx4, Mdlvx4, Tdlvx4, Aelvx4, Helvx4, Oelvx4, Velvx4, Cflvx4, Jflvx4, Qflvx4;
wire Xflvx4, Eglvx4, Lglvx4, Sglvx4, Zglvx4, Ghlvx4, Nhlvx4, Uhlvx4, Bilvx4, Iilvx4;
wire Pilvx4, Wilvx4, Djlvx4, Kjlvx4, Rjlvx4, Yjlvx4, Fklvx4, Mklvx4, Tklvx4, Allvx4;
wire Hllvx4, Ollvx4, Vllvx4, Cmlvx4, Jmlvx4, Qmlvx4, Xmlvx4, Enlvx4, Lnlvx4, Snlvx4;
wire Znlvx4, Golvx4, Nolvx4, Uolvx4, Bplvx4, Iplvx4, Pplvx4, Wplvx4, Dqlvx4, Kqlvx4;
wire Rqlvx4, Yqlvx4, Frlvx4, Mrlvx4, Trlvx4, Aslvx4, Hslvx4, Oslvx4, Vslvx4, Ctlvx4;
wire Jtlvx4, Qtlvx4, Xtlvx4, Eulvx4, Lulvx4, Sulvx4, Zulvx4, Gvlvx4, Nvlvx4, Uvlvx4;
wire Bwlvx4, Iwlvx4, Pwlvx4, Wwlvx4, Dxlvx4, Kxlvx4, Rxlvx4, Yxlvx4, Fylvx4, Mylvx4;
wire Tylvx4, Azlvx4, Hzlvx4, Ozlvx4, Vzlvx4, C0mvx4, J0mvx4, Q0mvx4, X0mvx4, E1mvx4;
wire L1mvx4, S1mvx4, Z1mvx4, G2mvx4, N2mvx4, U2mvx4, B3mvx4, I3mvx4, P3mvx4, W3mvx4;
wire D4mvx4, K4mvx4, R4mvx4, Y4mvx4, F5mvx4, M5mvx4, T5mvx4, A6mvx4, H6mvx4, O6mvx4;
wire V6mvx4, C7mvx4, J7mvx4, Q7mvx4, X7mvx4, E8mvx4, L8mvx4, S8mvx4, Z8mvx4, G9mvx4;
wire N9mvx4, U9mvx4, Bamvx4, Iamvx4, Pamvx4, Wamvx4, Dbmvx4, Kbmvx4, Rbmvx4, Ybmvx4;
wire Fcmvx4, Mcmvx4, Tcmvx4, Admvx4, Hdmvx4, Odmvx4, Vdmvx4, Cemvx4, Jemvx4, Qemvx4;
wire Xemvx4, Efmvx4, Lfmvx4, Sfmvx4, Zfmvx4, Ggmvx4, Ngmvx4, Ugmvx4, Bhmvx4, Ihmvx4;
wire Phmvx4, Whmvx4, Dimvx4, Kimvx4, Rimvx4, Yimvx4, Fjmvx4, Mjmvx4, Tjmvx4, Akmvx4;
wire Hkmvx4, Okmvx4, Vkmvx4, Clmvx4, Jlmvx4, Qlmvx4, Xlmvx4, Emmvx4, Lmmvx4, Smmvx4;
wire Zmmvx4, Gnmvx4, Nnmvx4, Unmvx4, Bomvx4, Iomvx4, Pomvx4, Womvx4, Dpmvx4, Kpmvx4;
wire Rpmvx4, Ypmvx4, Fqmvx4, Mqmvx4, Tqmvx4, Armvx4, Hrmvx4, Ormvx4, Vrmvx4, Csmvx4;
wire Jsmvx4, Qsmvx4, Xsmvx4, Etmvx4, Ltmvx4, Stmvx4, Ztmvx4, Gumvx4, Numvx4, Uumvx4;
wire Bvmvx4, Ivmvx4, Pvmvx4, Wvmvx4, Dwmvx4, Kwmvx4, Rwmvx4, Ywmvx4, Fxmvx4, Mxmvx4;
wire Txmvx4, Aymvx4, Hymvx4, Oymvx4, Vymvx4, Czmvx4, Jzmvx4, Qzmvx4, Xzmvx4, E0nvx4;
wire L0nvx4, S0nvx4, Z0nvx4, G1nvx4, N1nvx4, U1nvx4, B2nvx4, I2nvx4, P2nvx4, W2nvx4;
wire D3nvx4, K3nvx4, R3nvx4, Y3nvx4, F4nvx4, M4nvx4, T4nvx4, A5nvx4, H5nvx4, O5nvx4;
wire V5nvx4, C6nvx4, J6nvx4, Q6nvx4, X6nvx4, E7nvx4, L7nvx4, S7nvx4, Z7nvx4, G8nvx4;
wire N8nvx4, U8nvx4, B9nvx4, I9nvx4, P9nvx4, W9nvx4, Danvx4, Kanvx4, Ranvx4, Yanvx4;
wire Fbnvx4, Mbnvx4, Tbnvx4, Acnvx4, Hcnvx4, Ocnvx4, Vcnvx4, Cdnvx4, Jdnvx4, Qdnvx4;
wire Xdnvx4, Eenvx4, Lenvx4, Senvx4, Zenvx4, Gfnvx4, Nfnvx4, Ufnvx4, Bgnvx4, Ignvx4;
wire Pgnvx4, Wgnvx4, Dhnvx4, Khnvx4, Rhnvx4, Yhnvx4, Finvx4, Minvx4, Tinvx4, Ajnvx4;
wire Hjnvx4, Ojnvx4, Vjnvx4, Cknvx4, Jknvx4, Qknvx4, Xknvx4, Elnvx4, Llnvx4, Slnvx4;
wire Zlnvx4, Gmnvx4, Nmnvx4, Umnvx4, Bnnvx4, Innvx4, Pnnvx4, Wnnvx4, Donvx4, Konvx4;
wire Ronvx4, Yonvx4, Fpnvx4, Mpnvx4, Tpnvx4, Aqnvx4, Hqnvx4, Oqnvx4, Vqnvx4, Crnvx4;
wire Jrnvx4, Qrnvx4, Xrnvx4, Esnvx4, Lsnvx4, Ssnvx4, Zsnvx4, Gtnvx4, Ntnvx4, Utnvx4;
wire Bunvx4, Iunvx4, Punvx4, Wunvx4, Dvnvx4, Kvnvx4, Rvnvx4, Yvnvx4, Fwnvx4, Mwnvx4;
wire Twnvx4, Axnvx4, Hxnvx4, Oxnvx4, Vxnvx4, Cynvx4, Jynvx4, Qynvx4, Xynvx4, Eznvx4;
wire Lznvx4, Sznvx4, Zznvx4, G0ovx4, N0ovx4, U0ovx4, B1ovx4, I1ovx4, P1ovx4, W1ovx4;
wire D2ovx4, K2ovx4, R2ovx4, Y2ovx4, F3ovx4, M3ovx4, T3ovx4, A4ovx4, H4ovx4, O4ovx4;
wire V4ovx4, C5ovx4, J5ovx4, Q5ovx4, X5ovx4, E6ovx4, L6ovx4, S6ovx4, Z6ovx4, G7ovx4;
wire N7ovx4, U7ovx4, B8ovx4, I8ovx4, P8ovx4, W8ovx4, D9ovx4, K9ovx4, R9ovx4, Y9ovx4;
wire Faovx4, Maovx4, Taovx4, Abovx4, Hbovx4, Obovx4, Vbovx4, Ccovx4, Jcovx4, Qcovx4;
wire Xcovx4, Edovx4, Ldovx4, Sdovx4, Zdovx4, Geovx4, Neovx4, Ueovx4, Bfovx4, Ifovx4;
wire Pfovx4, Wfovx4, Dgovx4, Kgovx4, Rgovx4, Ygovx4, Fhovx4, Mhovx4, Thovx4, Aiovx4;
wire Hiovx4, Oiovx4, Viovx4, Cjovx4, Jjovx4, Qjovx4, Xjovx4, Ekovx4, Lkovx4, Skovx4;
wire Zkovx4, Glovx4, Nlovx4, Ulovx4, Bmovx4, Imovx4, Pmovx4, Wmovx4, Dnovx4, Knovx4;
wire Rnovx4, Ynovx4, Foovx4, Moovx4, Toovx4, Apovx4, Hpovx4, Opovx4, Vpovx4, Cqovx4;
wire Jqovx4, Qqovx4, Xqovx4, Erovx4, Lrovx4, Srovx4, Zrovx4, Gsovx4, Nsovx4, Usovx4;
wire Btovx4, Itovx4, Ptovx4, Wtovx4, Duovx4, Kuovx4, Ruovx4, Yuovx4, Fvovx4, Mvovx4;
wire Tvovx4, Awovx4, Hwovx4, Owovx4, Vwovx4, Cxovx4, Jxovx4, Qxovx4, Xxovx4, Eyovx4;
wire Lyovx4, Syovx4, Zyovx4, Gzovx4, Nzovx4, Uzovx4, B0pvx4, I0pvx4, P0pvx4, W0pvx4;
wire D1pvx4, K1pvx4, R1pvx4, Y1pvx4, F2pvx4, M2pvx4, T2pvx4, A3pvx4, H3pvx4, O3pvx4;
wire V3pvx4, C4pvx4, J4pvx4, Q4pvx4, X4pvx4, E5pvx4, L5pvx4, S5pvx4, Z5pvx4, G6pvx4;
wire N6pvx4, U6pvx4, B7pvx4, I7pvx4, P7pvx4, W7pvx4, D8pvx4, K8pvx4, R8pvx4, Y8pvx4;
wire F9pvx4, M9pvx4, T9pvx4, Aapvx4, Hapvx4, Oapvx4, Vapvx4, Cbpvx4, Jbpvx4, Qbpvx4;
wire Xbpvx4, Ecpvx4, Lcpvx4, Scpvx4, Zcpvx4, Gdpvx4, Ndpvx4, Udpvx4, Bepvx4, Iepvx4;
wire Pepvx4, Wepvx4, Dfpvx4, Kfpvx4, Rfpvx4, Yfpvx4, Fgpvx4, Mgpvx4, Tgpvx4, Ahpvx4;
wire Hhpvx4, Ohpvx4, Vhpvx4, Cipvx4, Jipvx4, Qipvx4, Xipvx4, Ejpvx4, Ljpvx4, Sjpvx4;
wire Zjpvx4, Gkpvx4, Nkpvx4, Ukpvx4, Blpvx4, Ilpvx4, Plpvx4, Wlpvx4, Dmpvx4, Kmpvx4;
wire Rmpvx4, Ympvx4, Fnpvx4, Mnpvx4, Tnpvx4, Aopvx4, Hopvx4, Oopvx4, Vopvx4, Cppvx4;
wire Jppvx4, Qppvx4, Xppvx4, Eqpvx4, Lqpvx4, Sqpvx4, Zqpvx4, Grpvx4, Nrpvx4, Urpvx4;
wire Bspvx4, Ispvx4, Pspvx4, Wspvx4, Dtpvx4, Ktpvx4, Rtpvx4, Ytpvx4, Fupvx4, Mupvx4;
wire Tupvx4, Avpvx4, Hvpvx4, Ovpvx4, Vvpvx4, Cwpvx4, Jwpvx4, Qwpvx4, Xwpvx4, Expvx4;
wire Lxpvx4, Sxpvx4, Zxpvx4, Gypvx4, Nypvx4, Uypvx4, Bzpvx4, Izpvx4, Pzpvx4, Wzpvx4;
wire D0qvx4, K0qvx4, R0qvx4, Y0qvx4, F1qvx4, M1qvx4, T1qvx4, A2qvx4, H2qvx4, O2qvx4;
wire V2qvx4, C3qvx4, J3qvx4, Q3qvx4, X3qvx4, E4qvx4, L4qvx4, S4qvx4, Z4qvx4, G5qvx4;
wire N5qvx4, U5qvx4, B6qvx4, I6qvx4, P6qvx4, W6qvx4, D7qvx4, K7qvx4, R7qvx4, Y7qvx4;
wire F8qvx4, M8qvx4, T8qvx4, A9qvx4, H9qvx4, O9qvx4, V9qvx4, Caqvx4, Jaqvx4, Qaqvx4;
wire Xaqvx4, Ebqvx4, Lbqvx4, Sbqvx4, Zbqvx4, Gcqvx4, Ncqvx4, Ucqvx4, Bdqvx4, Idqvx4;
wire Pdqvx4, Wdqvx4, Deqvx4, Keqvx4, Reqvx4, Yeqvx4, Ffqvx4, Mfqvx4, Tfqvx4, Agqvx4;
wire Hgqvx4, Ogqvx4, Vgqvx4, Chqvx4, Jhqvx4, Qhqvx4, Xhqvx4, Eiqvx4, Liqvx4, Siqvx4;
wire Ziqvx4, Gjqvx4, Njqvx4, Ujqvx4, Bkqvx4, Ikqvx4, Pkqvx4, Wkqvx4, Dlqvx4, Klqvx4;
wire Rlqvx4, Ylqvx4, Fmqvx4, Mmqvx4, Tmqvx4, Anqvx4, Hnqvx4, Onqvx4, Vnqvx4, Coqvx4;
wire Joqvx4, Qoqvx4, Xoqvx4, Epqvx4, Lpqvx4, Spqvx4, Zpqvx4, Gqqvx4, Nqqvx4, Uqqvx4;
wire Brqvx4, Irqvx4, Prqvx4, Wrqvx4, Dsqvx4, Ksqvx4, Rsqvx4, Ysqvx4, Ftqvx4, Mtqvx4;
wire Ttqvx4, Auqvx4, Huqvx4, Ouqvx4, Vuqvx4, Cvqvx4, Jvqvx4, Qvqvx4, Xvqvx4, Ewqvx4;
wire Lwqvx4, Swqvx4, Zwqvx4, Gxqvx4, Nxqvx4, Uxqvx4, Byqvx4, Iyqvx4, Pyqvx4, Wyqvx4;
wire Dzqvx4, Kzqvx4, Rzqvx4, Yzqvx4, F0rvx4, M0rvx4, T0rvx4, A1rvx4, H1rvx4, O1rvx4;
wire V1rvx4, C2rvx4, J2rvx4, Q2rvx4, X2rvx4, E3rvx4, L3rvx4, S3rvx4, Z3rvx4, G4rvx4;
wire N4rvx4, U4rvx4, B5rvx4, I5rvx4, P5rvx4, W5rvx4, D6rvx4, K6rvx4, R6rvx4, Y6rvx4;
wire F7rvx4, M7rvx4, T7rvx4, A8rvx4, H8rvx4, O8rvx4, V8rvx4, C9rvx4, J9rvx4, Q9rvx4;
wire X9rvx4, Earvx4, Larvx4, Sarvx4, Zarvx4, Gbrvx4, Nbrvx4, Ubrvx4, Bcrvx4, Icrvx4;
wire Pcrvx4, Wcrvx4, Ddrvx4, Kdrvx4, Rdrvx4, Ydrvx4, Fervx4, Mervx4, Tervx4, Afrvx4;
wire Hfrvx4, Ofrvx4, Vfrvx4, Cgrvx4, Jgrvx4, Qgrvx4, Xgrvx4, Ehrvx4, Lhrvx4, Shrvx4;
wire Zhrvx4, Girvx4, Nirvx4, Uirvx4, Bjrvx4, Ijrvx4, Pjrvx4, Wjrvx4, Dkrvx4, Kkrvx4;
wire Rkrvx4, Ykrvx4, Flrvx4, Mlrvx4, Tlrvx4, Amrvx4, Hmrvx4, Omrvx4, Vmrvx4, Cnrvx4;
wire Jnrvx4, Qnrvx4, Xnrvx4, Eorvx4, Lorvx4, Sorvx4, Zorvx4, Gprvx4, Nprvx4, Uprvx4;
wire Bqrvx4, Iqrvx4, Pqrvx4, Wqrvx4, Drrvx4, Krrvx4, Rrrvx4, Yrrvx4, Fsrvx4, Msrvx4;
wire Tsrvx4, Atrvx4, Htrvx4, Otrvx4, Vtrvx4, Curvx4, Jurvx4, Qurvx4, Xurvx4, Evrvx4;
wire Lvrvx4, Svrvx4, Zvrvx4, Gwrvx4, Nwrvx4, Uwrvx4, Bxrvx4, Ixrvx4, Pxrvx4, Wxrvx4;
wire Dyrvx4, Kyrvx4, Ryrvx4, Yyrvx4, Fzrvx4, Mzrvx4, Tzrvx4, A0svx4, H0svx4, O0svx4;
wire V0svx4, C1svx4, J1svx4, Q1svx4, X1svx4, E2svx4, L2svx4, S2svx4, Z2svx4, G3svx4;
wire N3svx4, U3svx4, B4svx4, I4svx4, P4svx4, W4svx4, D5svx4, K5svx4, R5svx4, Y5svx4;
wire F6svx4, M6svx4, T6svx4, A7svx4, H7svx4, O7svx4, V7svx4, C8svx4, J8svx4, Q8svx4;
wire X8svx4, E9svx4, L9svx4, S9svx4, Z9svx4, Gasvx4, Nasvx4, Uasvx4, Bbsvx4, Ibsvx4;
wire Pbsvx4, Wbsvx4, Dcsvx4, Kcsvx4, Rcsvx4, Ycsvx4, Fdsvx4, Mdsvx4, Tdsvx4, Aesvx4;
wire Hesvx4, Oesvx4, Vesvx4, Cfsvx4, Jfsvx4, Qfsvx4, Xfsvx4, Egsvx4, Lgsvx4, Sgsvx4;
wire Zgsvx4, Ghsvx4, Nhsvx4, Uhsvx4, Bisvx4, Iisvx4, Pisvx4, Wisvx4, Djsvx4, Kjsvx4;
wire Rjsvx4, Yjsvx4, Fksvx4, Mksvx4, Tksvx4, Alsvx4, Hlsvx4, Olsvx4, Vlsvx4, Cmsvx4;
wire Jmsvx4, Qmsvx4, Xmsvx4, Ensvx4, Lnsvx4, Snsvx4, Znsvx4, Gosvx4, Nosvx4, Uosvx4;
wire Bpsvx4, Ipsvx4, Ppsvx4, Wpsvx4, Dqsvx4, Kqsvx4, Rqsvx4, Yqsvx4, Frsvx4, Mrsvx4;
wire Trsvx4, Assvx4, Hssvx4, Ossvx4, Vssvx4, Ctsvx4, Jtsvx4, Qtsvx4, Xtsvx4, Eusvx4;
wire Lusvx4, Susvx4, Zusvx4, Gvsvx4, Nvsvx4, Uvsvx4, Bwsvx4, Iwsvx4, Pwsvx4, Wwsvx4;
wire Dxsvx4, Kxsvx4, Rxsvx4, Yxsvx4, Fysvx4, Mysvx4, Tysvx4, Azsvx4, Hzsvx4, Ozsvx4;
wire Vzsvx4, C0tvx4, J0tvx4, Q0tvx4, X0tvx4, E1tvx4, L1tvx4, S1tvx4, Z1tvx4, G2tvx4;
wire N2tvx4, U2tvx4, B3tvx4, I3tvx4, P3tvx4, W3tvx4, D4tvx4, K4tvx4, R4tvx4, Y4tvx4;
wire F5tvx4, M5tvx4, T5tvx4, A6tvx4, H6tvx4, O6tvx4, V6tvx4, C7tvx4, J7tvx4, Q7tvx4;
wire X7tvx4, E8tvx4, L8tvx4, S8tvx4, Z8tvx4, G9tvx4, N9tvx4, U9tvx4, Batvx4, Iatvx4;
wire Patvx4, Watvx4, Dbtvx4, Kbtvx4, Rbtvx4, Ybtvx4, Fctvx4, Mctvx4, Tctvx4, Adtvx4;
wire Hdtvx4, Odtvx4, Vdtvx4, Cetvx4, Jetvx4, Qetvx4, Xetvx4, Eftvx4, Lftvx4, Sftvx4;
wire Zftvx4, Ggtvx4, Ngtvx4, Ugtvx4, Bhtvx4, Ihtvx4, Phtvx4, Whtvx4, Ditvx4, Kitvx4;
wire Ritvx4, Yitvx4, Fjtvx4, Mjtvx4, Tjtvx4, Aktvx4, Hktvx4, Oktvx4, Vktvx4, Cltvx4;
wire Jltvx4, Qltvx4, Xltvx4, Emtvx4, Lmtvx4, Smtvx4, Zmtvx4, Gntvx4, Nntvx4, Untvx4;
wire Botvx4, Iotvx4, Potvx4, Wotvx4, Dptvx4, Kptvx4, Rptvx4, Yptvx4, Fqtvx4, Mqtvx4;
wire Tqtvx4, Artvx4, Hrtvx4, Ortvx4, Vrtvx4, Cstvx4, Jstvx4, Qstvx4, Xstvx4, Ettvx4;
wire Lttvx4, Sttvx4, Zttvx4, Gutvx4, Nutvx4, Uutvx4, Bvtvx4, Ivtvx4, Pvtvx4, Wvtvx4;
wire Dwtvx4, Kwtvx4, Rwtvx4, Ywtvx4, Fxtvx4, Mxtvx4, Txtvx4, Aytvx4, Hytvx4, Oytvx4;
wire Vytvx4, Cztvx4, Jztvx4, Qztvx4, Xztvx4, E0uvx4, L0uvx4, S0uvx4, Z0uvx4, G1uvx4;
wire N1uvx4, U1uvx4, B2uvx4, I2uvx4, P2uvx4, W2uvx4, D3uvx4, K3uvx4, R3uvx4, Y3uvx4;
wire F4uvx4, M4uvx4, T4uvx4, A5uvx4, H5uvx4, O5uvx4, V5uvx4, C6uvx4, J6uvx4, Q6uvx4;
wire X6uvx4, E7uvx4, L7uvx4, S7uvx4, Z7uvx4, G8uvx4, N8uvx4, U8uvx4, B9uvx4, I9uvx4;
wire P9uvx4, W9uvx4, Dauvx4, Kauvx4, Rauvx4, Yauvx4, Fbuvx4, Mbuvx4, Tbuvx4, Acuvx4;
wire Hcuvx4, Ocuvx4, Vcuvx4, Cduvx4, Jduvx4, Qduvx4, Xduvx4, Eeuvx4, Leuvx4, Seuvx4;
wire Zeuvx4, Gfuvx4, Nfuvx4, Ufuvx4, Bguvx4, Iguvx4, Pguvx4, Wguvx4, Dhuvx4, Khuvx4;
wire Rhuvx4, Yhuvx4, Fiuvx4, Miuvx4, Tiuvx4, Ajuvx4, Hjuvx4, Ojuvx4, Vjuvx4, Ckuvx4;
wire Jkuvx4, Qkuvx4, Xkuvx4, Eluvx4, Lluvx4, Sluvx4, Zluvx4, Gmuvx4, Nmuvx4, Umuvx4;
wire Bnuvx4, Inuvx4, Pnuvx4, Wnuvx4, Douvx4, Kouvx4, Rouvx4, Youvx4, Fpuvx4, Mpuvx4;
wire Tpuvx4, Aquvx4, Hquvx4, Oquvx4, Vquvx4, Cruvx4, Jruvx4, Qruvx4, Xruvx4, Esuvx4;
wire Lsuvx4, Ssuvx4, Zsuvx4, Gtuvx4, Ntuvx4, Utuvx4, Buuvx4, Iuuvx4, Puuvx4, Wuuvx4;
wire Dvuvx4, Kvuvx4, Rvuvx4, Yvuvx4, Fwuvx4, Mwuvx4, Twuvx4, Axuvx4, Hxuvx4, Oxuvx4;
wire Vxuvx4, Cyuvx4, Jyuvx4, Qyuvx4, Xyuvx4, Ezuvx4, Lzuvx4, Szuvx4, Zzuvx4, G0vvx4;
wire N0vvx4, U0vvx4, B1vvx4, I1vvx4, P1vvx4, W1vvx4, D2vvx4, K2vvx4, R2vvx4, Y2vvx4;
wire F3vvx4, M3vvx4, T3vvx4, A4vvx4, H4vvx4, O4vvx4, V4vvx4, C5vvx4, J5vvx4, Q5vvx4;
wire X5vvx4, E6vvx4, L6vvx4, S6vvx4, Z6vvx4, G7vvx4, N7vvx4, U7vvx4, B8vvx4, I8vvx4;
wire P8vvx4, W8vvx4, D9vvx4, K9vvx4, R9vvx4, Y9vvx4, Favvx4, Mavvx4, Tavvx4, Abvvx4;
wire Hbvvx4, Obvvx4, Vbvvx4, Ccvvx4, Jcvvx4, Qcvvx4, Xcvvx4, Edvvx4, Ldvvx4, Sdvvx4;
wire Zdvvx4, Gevvx4, Nevvx4, Uevvx4, Bfvvx4, Ifvvx4, Pfvvx4, Wfvvx4, Dgvvx4, Kgvvx4;
wire Rgvvx4, Ygvvx4, Fhvvx4, Mhvvx4, Thvvx4, Aivvx4, Hivvx4, Oivvx4, Vivvx4, Cjvvx4;
wire Jjvvx4, Qjvvx4, Xjvvx4, Ekvvx4, Lkvvx4, Skvvx4, Zkvvx4, Glvvx4, Nlvvx4, Ulvvx4;
wire Bmvvx4, Imvvx4, Pmvvx4, Wmvvx4, Dnvvx4, Knvvx4, Rnvvx4, Ynvvx4, Fovvx4, Movvx4;
wire Tovvx4, Apvvx4, Hpvvx4, Opvvx4, Vpvvx4, Cqvvx4, Jqvvx4, Qqvvx4, Xqvvx4, Ervvx4;
wire Lrvvx4, Srvvx4, Zrvvx4, Gsvvx4, Nsvvx4, Usvvx4, Btvvx4, Itvvx4, Ptvvx4, Wtvvx4;
wire Duvvx4, Kuvvx4, Ruvvx4, Yuvvx4, Fvvvx4, Mvvvx4, Tvvvx4, Awvvx4, Hwvvx4, Owvvx4;
wire Vwvvx4, Cxvvx4, Jxvvx4, Qxvvx4, Xxvvx4, Eyvvx4, Lyvvx4, Syvvx4, Zyvvx4, Gzvvx4;
wire Nzvvx4, Uzvvx4, B0wvx4, I0wvx4, P0wvx4, W0wvx4, D1wvx4, K1wvx4, R1wvx4, Y1wvx4;
wire F2wvx4, M2wvx4, T2wvx4, A3wvx4, H3wvx4, O3wvx4, V3wvx4, C4wvx4, J4wvx4, Q4wvx4;
wire X4wvx4, E5wvx4, L5wvx4, S5wvx4, Z5wvx4, G6wvx4, N6wvx4, U6wvx4, B7wvx4, I7wvx4;
wire P7wvx4, W7wvx4, D8wvx4, K8wvx4, R8wvx4, Y8wvx4, F9wvx4, M9wvx4, T9wvx4, Aawvx4;
wire Hawvx4, Oawvx4, Vawvx4, Cbwvx4, Jbwvx4, Qbwvx4, Xbwvx4, Ecwvx4, Lcwvx4, Scwvx4;
wire Zcwvx4, Gdwvx4, Ndwvx4, Udwvx4, Bewvx4, Iewvx4, Pewvx4, Wewvx4, Dfwvx4, Kfwvx4;
wire Rfwvx4, Yfwvx4, Fgwvx4, Mgwvx4, Tgwvx4, Ahwvx4, Hhwvx4, Ohwvx4, Vhwvx4, Ciwvx4;
wire Jiwvx4, Qiwvx4, Xiwvx4, Ejwvx4, Ljwvx4, Sjwvx4, Zjwvx4, Gkwvx4, Nkwvx4, Ukwvx4;
wire Blwvx4, Ilwvx4, Plwvx4, Wlwvx4, Dmwvx4, Kmwvx4, Rmwvx4, Ymwvx4, Fnwvx4, Mnwvx4;
wire Tnwvx4, Aowvx4, Howvx4, Oowvx4, Vowvx4, Cpwvx4, Jpwvx4, Qpwvx4, Xpwvx4, Eqwvx4;
wire Lqwvx4, Sqwvx4, Zqwvx4, Grwvx4, Nrwvx4, Urwvx4, Bswvx4, Iswvx4, Pswvx4, Wswvx4;
wire Dtwvx4, Ktwvx4, Rtwvx4, Ytwvx4, Fuwvx4, Muwvx4, Tuwvx4, Avwvx4, Hvwvx4, Ovwvx4;
wire Vvwvx4, Cwwvx4, Jwwvx4, Qwwvx4, Xwwvx4, Exwvx4, Lxwvx4, Sxwvx4, Zxwvx4, Gywvx4;
wire Nywvx4, Uywvx4, Bzwvx4, Izwvx4, Pzwvx4, Wzwvx4, D0xvx4, K0xvx4, R0xvx4, Y0xvx4;
wire F1xvx4, M1xvx4, T1xvx4, A2xvx4, H2xvx4, O2xvx4, V2xvx4, C3xvx4, J3xvx4, Q3xvx4;
wire X3xvx4, E4xvx4, L4xvx4, S4xvx4, Z4xvx4, G5xvx4, N5xvx4, U5xvx4, B6xvx4, I6xvx4;
wire P6xvx4, W6xvx4, D7xvx4, K7xvx4, R7xvx4, Y7xvx4, F8xvx4, M8xvx4, T8xvx4, A9xvx4;
wire H9xvx4, O9xvx4, V9xvx4, Caxvx4, Jaxvx4, Qaxvx4, Xaxvx4, Ebxvx4, Lbxvx4, Sbxvx4;
wire Zbxvx4, Gcxvx4, Ncxvx4, Ucxvx4, Bdxvx4, Idxvx4, Pdxvx4, Wdxvx4, Dexvx4, Kexvx4;
wire Rexvx4, Yexvx4, Ffxvx4, Mfxvx4, Tfxvx4, Agxvx4, Hgxvx4, Ogxvx4, Vgxvx4, Chxvx4;
wire Jhxvx4, Qhxvx4, Xhxvx4, Eixvx4, Lixvx4, Sixvx4, Zixvx4, Gjxvx4, Njxvx4, Ujxvx4;
wire Bkxvx4, Ikxvx4, Pkxvx4, Wkxvx4, Dlxvx4, Klxvx4, Rlxvx4, Ylxvx4, Fmxvx4, Mmxvx4;
wire Tmxvx4, Anxvx4, Hnxvx4, Onxvx4, Vnxvx4, Coxvx4, Joxvx4, Qoxvx4, Xoxvx4, Epxvx4;
wire Lpxvx4, Spxvx4, Zpxvx4, Gqxvx4, Nqxvx4, Uqxvx4, Brxvx4, Irxvx4, Prxvx4, Wrxvx4;
wire Dsxvx4, Ksxvx4, Rsxvx4, Ysxvx4, Ftxvx4, Mtxvx4, Ttxvx4, Auxvx4, Huxvx4, Ouxvx4;
wire Vuxvx4, Cvxvx4, Jvxvx4, Qvxvx4, Xvxvx4, Ewxvx4, Lwxvx4, Swxvx4, Zwxvx4, Gxxvx4;
wire Nxxvx4, Uxxvx4, Byxvx4, Iyxvx4, Pyxvx4, Wyxvx4, Dzxvx4, Kzxvx4, Rzxvx4, Yzxvx4;
wire F0yvx4, M0yvx4, T0yvx4, A1yvx4, H1yvx4, O1yvx4, V1yvx4, C2yvx4, J2yvx4, Q2yvx4;
wire X2yvx4, E3yvx4, L3yvx4, S3yvx4, Z3yvx4, G4yvx4, N4yvx4, U4yvx4, B5yvx4, I5yvx4;
wire P5yvx4, W5yvx4, D6yvx4, K6yvx4, R6yvx4, Y6yvx4, F7yvx4, M7yvx4, T7yvx4, A8yvx4;
wire H8yvx4, O8yvx4, V8yvx4, C9yvx4, J9yvx4, Q9yvx4, X9yvx4, Eayvx4, Layvx4, Sayvx4;
wire Zayvx4, Gbyvx4, Nbyvx4, Ubyvx4, Bcyvx4, Icyvx4, Pcyvx4, Wcyvx4, Ddyvx4, Kdyvx4;
wire Rdyvx4, Ydyvx4, Feyvx4, Meyvx4, Teyvx4, Afyvx4, Hfyvx4, Ofyvx4, Vfyvx4, Cgyvx4;
wire Jgyvx4, Qgyvx4, Xgyvx4, Ehyvx4, Lhyvx4, Shyvx4, Zhyvx4, Giyvx4, Niyvx4, Uiyvx4;
wire Bjyvx4, Ijyvx4, Pjyvx4, Wjyvx4, Dkyvx4, Kkyvx4, Rkyvx4, Ykyvx4, Flyvx4, Mlyvx4;
wire Tlyvx4, Amyvx4, Hmyvx4, Omyvx4, Vmyvx4, Cnyvx4, Jnyvx4, Qnyvx4, Xnyvx4, Eoyvx4;
wire Loyvx4, Soyvx4, Zoyvx4, Gpyvx4, Npyvx4, Upyvx4, Bqyvx4, Iqyvx4, Pqyvx4, Wqyvx4;
wire Dryvx4, Kryvx4, Rryvx4, Yryvx4, Fsyvx4, Msyvx4, Tsyvx4, Atyvx4, Htyvx4, Otyvx4;
wire Vtyvx4, Cuyvx4, Juyvx4, Quyvx4, Xuyvx4, Evyvx4, Lvyvx4, Svyvx4, Zvyvx4, Gwyvx4;
wire Nwyvx4, Uwyvx4, Bxyvx4, Ixyvx4, Pxyvx4, Wxyvx4, Dyyvx4, Kyyvx4, Ryyvx4, Yyyvx4;
wire Fzyvx4, Mzyvx4, Tzyvx4, A0zvx4, H0zvx4, O0zvx4, V0zvx4, C1zvx4, J1zvx4, Q1zvx4;
wire X1zvx4, E2zvx4, L2zvx4, S2zvx4, Z2zvx4, G3zvx4, N3zvx4, U3zvx4, B4zvx4, I4zvx4;
wire P4zvx4, W4zvx4, D5zvx4, K5zvx4, R5zvx4, Y5zvx4, F6zvx4, M6zvx4, T6zvx4, A7zvx4;
wire H7zvx4, O7zvx4, V7zvx4, C8zvx4, J8zvx4, Q8zvx4, X8zvx4, E9zvx4, L9zvx4, S9zvx4;
wire Z9zvx4, Gazvx4, Nazvx4, Uazvx4, Bbzvx4, Ibzvx4, Pbzvx4, Wbzvx4, Dczvx4, Kczvx4;
wire Rczvx4, Yczvx4, Fdzvx4, Mdzvx4, Tdzvx4, Aezvx4, Hezvx4, Oezvx4, Vezvx4, Cfzvx4;
wire Jfzvx4, Qfzvx4, Xfzvx4, Egzvx4, Lgzvx4, Sgzvx4, Zgzvx4, Ghzvx4, Nhzvx4, Uhzvx4;
wire Bizvx4, Iizvx4, Pizvx4, Wizvx4, Djzvx4, Kjzvx4, Rjzvx4, Yjzvx4, Fkzvx4, Mkzvx4;
wire Tkzvx4, Alzvx4, Hlzvx4, Olzvx4, Vlzvx4, Cmzvx4, Jmzvx4, Qmzvx4, Xmzvx4, Enzvx4;
wire Lnzvx4, Snzvx4, Znzvx4, Gozvx4, Nozvx4, Uozvx4, Bpzvx4, Ipzvx4, Ppzvx4, Wpzvx4;
wire Dqzvx4, Kqzvx4, Rqzvx4, Yqzvx4, Frzvx4, Mrzvx4, Trzvx4, Aszvx4, Hszvx4, Oszvx4;
wire Vszvx4, Ctzvx4, Jtzvx4, Qtzvx4, Xtzvx4, Euzvx4, Luzvx4, Suzvx4, Zuzvx4, Gvzvx4;
wire Nvzvx4, Uvzvx4, Bwzvx4, Iwzvx4, Pwzvx4, Wwzvx4, Dxzvx4, Kxzvx4, Rxzvx4, Yxzvx4;
wire Fyzvx4, Myzvx4, Tyzvx4, Azzvx4, Hzzvx4, Ozzvx4, Vzzvx4, C00wx4, J00wx4, Q00wx4;
wire X00wx4, E10wx4, L10wx4, S10wx4, Z10wx4, G20wx4, N20wx4, U20wx4, B30wx4, I30wx4;
wire P30wx4, W30wx4, D40wx4, K40wx4, R40wx4, Y40wx4, F50wx4, M50wx4, T50wx4, A60wx4;
wire H60wx4, O60wx4, V60wx4, C70wx4, J70wx4, Q70wx4, X70wx4, E80wx4, L80wx4, S80wx4;
wire Z80wx4, G90wx4, N90wx4, U90wx4, Ba0wx4, Ia0wx4, Pa0wx4, Wa0wx4, Db0wx4, Kb0wx4;
wire Rb0wx4, Yb0wx4, Fc0wx4, Mc0wx4, Tc0wx4, Ad0wx4, Hd0wx4, Od0wx4, Vd0wx4, Ce0wx4;
wire Je0wx4, Qe0wx4, Xe0wx4, Ef0wx4, Lf0wx4, Sf0wx4, Zf0wx4, Gg0wx4, Ng0wx4, Ug0wx4;
wire Bh0wx4, Ih0wx4, Ph0wx4, Wh0wx4, Di0wx4, Ki0wx4, Ri0wx4, Yi0wx4, Fj0wx4, Mj0wx4;
wire Tj0wx4, Ak0wx4, Hk0wx4, Ok0wx4, Vk0wx4, Cl0wx4, Jl0wx4, Ql0wx4, Xl0wx4, Em0wx4;
wire Lm0wx4, Sm0wx4, Zm0wx4, Gn0wx4, Nn0wx4, Un0wx4, Bo0wx4, Io0wx4, Po0wx4, Wo0wx4;
wire Dp0wx4, Kp0wx4, Rp0wx4, Yp0wx4, Fq0wx4, Mq0wx4, Tq0wx4, Ar0wx4, Hr0wx4, Or0wx4;
wire Vr0wx4, Cs0wx4, Js0wx4, Qs0wx4, Xs0wx4, Et0wx4, Lt0wx4, St0wx4, Zt0wx4, Gu0wx4;
wire Nu0wx4, Uu0wx4, Bv0wx4, Iv0wx4, Pv0wx4, Wv0wx4, Dw0wx4, Kw0wx4, Rw0wx4, Yw0wx4;
wire Fx0wx4, Mx0wx4, Tx0wx4, Ay0wx4, Hy0wx4, Oy0wx4, Vy0wx4, Cz0wx4, Jz0wx4, Qz0wx4;
wire Xz0wx4, E01wx4, L01wx4, S01wx4, Z01wx4, G11wx4, N11wx4, U11wx4, B21wx4, I21wx4;
wire P21wx4, W21wx4, D31wx4, K31wx4, R31wx4, Y31wx4, F41wx4, M41wx4, T41wx4, A51wx4;
wire H51wx4, O51wx4, V51wx4, C61wx4, J61wx4, Q61wx4, X61wx4, E71wx4, L71wx4, S71wx4;
wire Z71wx4, G81wx4, N81wx4, U81wx4, B91wx4, I91wx4, P91wx4, W91wx4, Da1wx4, Ka1wx4;
wire Ra1wx4, Ya1wx4, Fb1wx4, Mb1wx4, Tb1wx4, Ac1wx4, Hc1wx4, Oc1wx4, Vc1wx4, Cd1wx4;
wire Jd1wx4, Qd1wx4, Xd1wx4, Ee1wx4, Le1wx4, Se1wx4, Ze1wx4, Gf1wx4, Nf1wx4, Uf1wx4;
wire Bg1wx4, Ig1wx4, Pg1wx4, Wg1wx4, Dh1wx4, Kh1wx4, Rh1wx4, Yh1wx4, Fi1wx4, Mi1wx4;
wire Ti1wx4, Aj1wx4, Hj1wx4, Oj1wx4, Vj1wx4, Ck1wx4, Jk1wx4, Qk1wx4, Xk1wx4, El1wx4;
wire Ll1wx4, Sl1wx4, Zl1wx4, Gm1wx4, Nm1wx4, Um1wx4, Bn1wx4, In1wx4, Pn1wx4, Wn1wx4;
wire Do1wx4, Ko1wx4, Ro1wx4, Yo1wx4, Fp1wx4, Mp1wx4, Tp1wx4, Aq1wx4, Hq1wx4, Oq1wx4;
wire Vq1wx4, Cr1wx4, Jr1wx4, Qr1wx4, Xr1wx4, Es1wx4, Ls1wx4, Ss1wx4, Zs1wx4, Gt1wx4;
wire Nt1wx4, Ut1wx4, Bu1wx4, Iu1wx4, Pu1wx4, Wu1wx4, Dv1wx4, Kv1wx4, Rv1wx4, Yv1wx4;
wire Fw1wx4, Mw1wx4, Tw1wx4, Ax1wx4, Hx1wx4, Ox1wx4, Vx1wx4, Cy1wx4, Jy1wx4, Qy1wx4;
wire Xy1wx4, Ez1wx4, Lz1wx4, Sz1wx4, Zz1wx4, G02wx4, N02wx4, U02wx4, B12wx4, I12wx4;
wire P12wx4, W12wx4, D22wx4, K22wx4, R22wx4, Y22wx4, F32wx4, M32wx4, T32wx4, A42wx4;
wire H42wx4, O42wx4, V42wx4, C52wx4, J52wx4, Q52wx4, X52wx4, E62wx4, L62wx4, S62wx4;
wire Z62wx4, G72wx4, N72wx4, U72wx4, B82wx4, I82wx4, P82wx4, W82wx4, D92wx4, K92wx4;
wire R92wx4, Y92wx4, Fa2wx4, Ma2wx4, Ta2wx4, Ab2wx4, Hb2wx4, Ob2wx4, Vb2wx4, Cc2wx4;
wire Jc2wx4, Qc2wx4, Xc2wx4, Ed2wx4, Ld2wx4, Sd2wx4, Zd2wx4, Ge2wx4, Ne2wx4, Ue2wx4;
wire Bf2wx4, If2wx4, Pf2wx4, Wf2wx4, Dg2wx4, Kg2wx4, Rg2wx4, Yg2wx4, Fh2wx4, Mh2wx4;
wire Th2wx4, Ai2wx4, Hi2wx4, Oi2wx4, Vi2wx4, Cj2wx4, Jj2wx4, Qj2wx4, Xj2wx4, Ek2wx4;
wire Lk2wx4, Sk2wx4, Zk2wx4, Gl2wx4, Nl2wx4, Ul2wx4, Bm2wx4, Im2wx4, Pm2wx4, Wm2wx4;
wire Dn2wx4, Kn2wx4, Rn2wx4, Yn2wx4, Fo2wx4, Mo2wx4, To2wx4, Ap2wx4, Hp2wx4, Op2wx4;
wire Vp2wx4, Cq2wx4, Jq2wx4, Qq2wx4, Xq2wx4, Er2wx4, Lr2wx4, Sr2wx4, Zr2wx4, Gs2wx4;
wire Ns2wx4, Us2wx4, Bt2wx4, It2wx4, Pt2wx4, Wt2wx4, Du2wx4, Ku2wx4, Ru2wx4, Yu2wx4;
wire Fv2wx4, Mv2wx4, Tv2wx4, Aw2wx4, Hw2wx4, Ow2wx4, Vw2wx4, Cx2wx4, Jx2wx4, Qx2wx4;
wire Xx2wx4, Ey2wx4, Ly2wx4, Sy2wx4, Zy2wx4, Gz2wx4, Nz2wx4, Uz2wx4, B03wx4, I03wx4;
wire P03wx4, W03wx4, D13wx4, K13wx4, R13wx4, Y13wx4, F23wx4, M23wx4, T23wx4, A33wx4;
wire H33wx4, O33wx4, V33wx4, C43wx4, J43wx4, Q43wx4, X43wx4, E53wx4, L53wx4, S53wx4;
wire Z53wx4, G63wx4, N63wx4, U63wx4, B73wx4, I73wx4, P73wx4, W73wx4, D83wx4, K83wx4;
wire R83wx4, Y83wx4, F93wx4, M93wx4, T93wx4, Aa3wx4, Ha3wx4, Oa3wx4, Va3wx4, Cb3wx4;
wire Jb3wx4, Qb3wx4, Xb3wx4, Ec3wx4, Lc3wx4, Sc3wx4, Zc3wx4, Gd3wx4, Nd3wx4, Ud3wx4;
wire Be3wx4, Ie3wx4, Pe3wx4, We3wx4, Df3wx4, Kf3wx4, Rf3wx4, Yf3wx4, Fg3wx4, Mg3wx4;
wire Tg3wx4, Ah3wx4, Hh3wx4, Oh3wx4, Vh3wx4, Ci3wx4, Ji3wx4, Qi3wx4, Xi3wx4, Ej3wx4;
wire Lj3wx4, Sj3wx4, Zj3wx4, Gk3wx4, Nk3wx4, Uk3wx4, Bl3wx4, Il3wx4, Pl3wx4, Wl3wx4;
wire Dm3wx4, Km3wx4, Rm3wx4, Ym3wx4, Fn3wx4, Mn3wx4, Tn3wx4, Ao3wx4, Ho3wx4, Oo3wx4;
wire Vo3wx4, Cp3wx4, Jp3wx4, Qp3wx4, Xp3wx4, Eq3wx4, Lq3wx4, Sq3wx4, Zq3wx4, Gr3wx4;
wire Nr3wx4, Ur3wx4, Bs3wx4, Is3wx4, Ps3wx4, Ws3wx4, Dt3wx4, Kt3wx4, Rt3wx4, Yt3wx4;
wire Fu3wx4, Mu3wx4, Tu3wx4, Av3wx4, Hv3wx4, Ov3wx4, Vv3wx4, Cw3wx4, Jw3wx4, Qw3wx4;
wire Xw3wx4, Ex3wx4, Lx3wx4, Sx3wx4, Zx3wx4, Gy3wx4, Ny3wx4, Uy3wx4, Bz3wx4, Iz3wx4;
wire Pz3wx4, Wz3wx4, D04wx4, K04wx4, R04wx4, Y04wx4, F14wx4, M14wx4, T14wx4, A24wx4;
wire H24wx4, O24wx4, V24wx4, C34wx4, J34wx4, Q34wx4, X34wx4, E44wx4, L44wx4, S44wx4;
wire Z44wx4, G54wx4, N54wx4, U54wx4, B64wx4, I64wx4, P64wx4, W64wx4, D74wx4, K74wx4;
wire R74wx4, Y74wx4, F84wx4, M84wx4, T84wx4, A94wx4, H94wx4, O94wx4, V94wx4, Ca4wx4;
wire Ja4wx4, Qa4wx4, Xa4wx4, Eb4wx4, Lb4wx4, Sb4wx4, Zb4wx4, Gc4wx4, Nc4wx4, Uc4wx4;
wire Bd4wx4, Id4wx4, Pd4wx4, Wd4wx4, De4wx4, Ke4wx4, Re4wx4, Ye4wx4, Ff4wx4, Mf4wx4;
wire Tf4wx4, Ag4wx4, Hg4wx4, Og4wx4, Vg4wx4, Ch4wx4, Jh4wx4, Qh4wx4, Xh4wx4, Ei4wx4;
wire Li4wx4, Si4wx4, Zi4wx4, Gj4wx4, Nj4wx4, Uj4wx4, Bk4wx4, Ik4wx4, Pk4wx4, Wk4wx4;
wire Dl4wx4, Kl4wx4, Rl4wx4, Yl4wx4, Fm4wx4, Mm4wx4, Tm4wx4, An4wx4, Hn4wx4, On4wx4;
wire Vn4wx4, Co4wx4, Jo4wx4, Qo4wx4, Xo4wx4, Ep4wx4, Lp4wx4, Sp4wx4, Zp4wx4, Gq4wx4;
wire Nq4wx4, Uq4wx4, Br4wx4, Ir4wx4, Pr4wx4, Wr4wx4, Ds4wx4, Ks4wx4, Rs4wx4, Ys4wx4;
wire Ft4wx4, Mt4wx4, Tt4wx4, Au4wx4, Hu4wx4, Ou4wx4, Vu4wx4, Cv4wx4, Jv4wx4, Qv4wx4;
wire Xv4wx4, Ew4wx4, Lw4wx4, Sw4wx4, Zw4wx4, Gx4wx4, Nx4wx4, Ux4wx4, By4wx4, Iy4wx4;
wire Py4wx4, Wy4wx4, Dz4wx4, Kz4wx4, Rz4wx4, Yz4wx4, F05wx4, M05wx4, T05wx4, A15wx4;
wire H15wx4, O15wx4, V15wx4, C25wx4, J25wx4, Q25wx4, X25wx4, E35wx4, L35wx4, S35wx4;
wire Z35wx4, G45wx4, N45wx4, U45wx4, B55wx4, I55wx4, P55wx4, W55wx4, D65wx4, K65wx4;
wire R65wx4, Y65wx4, F75wx4, M75wx4, T75wx4, A85wx4, H85wx4, O85wx4, V85wx4, C95wx4;
wire J95wx4, Q95wx4, X95wx4, Ea5wx4, La5wx4, Sa5wx4, Za5wx4, Gb5wx4, Nb5wx4, Ub5wx4;
wire Bc5wx4, Ic5wx4, Pc5wx4, Wc5wx4, Dd5wx4, Kd5wx4, Rd5wx4, Yd5wx4, Fe5wx4, Me5wx4;
wire Te5wx4, Af5wx4, Hf5wx4, Of5wx4, Vf5wx4, Cg5wx4, Jg5wx4, Qg5wx4, Xg5wx4, Eh5wx4;
wire Lh5wx4, Sh5wx4, Zh5wx4, Gi5wx4, Ni5wx4, Ui5wx4, Bj5wx4, Ij5wx4, Pj5wx4, Wj5wx4;
wire Dk5wx4, Kk5wx4, Rk5wx4, Yk5wx4, Fl5wx4, Ml5wx4, Tl5wx4, Am5wx4, Hm5wx4, Om5wx4;
wire Vm5wx4, Cn5wx4, Jn5wx4, Qn5wx4, Xn5wx4, Eo5wx4, Lo5wx4, So5wx4, Zo5wx4, Gp5wx4;
wire Np5wx4, Up5wx4, Bq5wx4, Iq5wx4, Pq5wx4, Wq5wx4, Dr5wx4, Kr5wx4, Rr5wx4, Yr5wx4;
wire Fs5wx4, Ms5wx4, Ts5wx4, At5wx4, Ht5wx4, Ot5wx4, Vt5wx4, Cu5wx4, Ju5wx4, Qu5wx4;
wire Xu5wx4, Ev5wx4, Lv5wx4, Sv5wx4, Zv5wx4, Gw5wx4, Nw5wx4, Uw5wx4, Bx5wx4, Ix5wx4;
wire Px5wx4, Wx5wx4, Dy5wx4, Ky5wx4, Ry5wx4, Yy5wx4, Fz5wx4, Mz5wx4, Tz5wx4, A06wx4;
wire H06wx4, O06wx4, V06wx4, C16wx4, J16wx4, Q16wx4, X16wx4, E26wx4, L26wx4, S26wx4;
wire Z26wx4, G36wx4, N36wx4, U36wx4, B46wx4, I46wx4, P46wx4, W46wx4, D56wx4, K56wx4;
wire R56wx4, Y56wx4, F66wx4, M66wx4, T66wx4, A76wx4, H76wx4, O76wx4, V76wx4, C86wx4;
wire J86wx4, Q86wx4, X86wx4, E96wx4, L96wx4, S96wx4, Z96wx4, Ga6wx4, Na6wx4, Ua6wx4;
wire Bb6wx4, Ib6wx4, Pb6wx4, Wb6wx4, Dc6wx4, Kc6wx4, Rc6wx4, Yc6wx4, Fd6wx4, Md6wx4;
wire Td6wx4, Ae6wx4, He6wx4, Oe6wx4, Ve6wx4, Cf6wx4, Jf6wx4, Qf6wx4, Xf6wx4, Eg6wx4;
wire Lg6wx4, Sg6wx4, Zg6wx4, Gh6wx4, Nh6wx4, Uh6wx4, Bi6wx4, Ii6wx4, Pi6wx4, Wi6wx4;
wire Dj6wx4, Kj6wx4, Rj6wx4, Yj6wx4, Fk6wx4, Mk6wx4, Tk6wx4, Al6wx4, Hl6wx4, Ol6wx4;
wire Vl6wx4, Cm6wx4, Jm6wx4, Qm6wx4, Xm6wx4, En6wx4, Ln6wx4, Sn6wx4, Zn6wx4, Go6wx4;
wire No6wx4, Uo6wx4, Bp6wx4, Ip6wx4, Pp6wx4, Wp6wx4, Dq6wx4, Kq6wx4, Rq6wx4, Yq6wx4;
wire Fr6wx4, Mr6wx4, Tr6wx4, As6wx4, Hs6wx4, Os6wx4, Vs6wx4, Ct6wx4, Jt6wx4, Qt6wx4;
wire Xt6wx4, Eu6wx4, Lu6wx4, Su6wx4, Zu6wx4, Gv6wx4, Nv6wx4, Uv6wx4, Bw6wx4, Iw6wx4;
wire Pw6wx4, Ww6wx4, Dx6wx4, Kx6wx4, Rx6wx4, Yx6wx4, Fy6wx4, My6wx4, Ty6wx4, Az6wx4;
wire Hz6wx4, Oz6wx4, Vz6wx4, C07wx4, J07wx4, Q07wx4, X07wx4, E17wx4, L17wx4, S17wx4;
wire Z17wx4, G27wx4, N27wx4, U27wx4, B37wx4, I37wx4, P37wx4, W37wx4, D47wx4, K47wx4;
wire R47wx4, Y47wx4, F57wx4, M57wx4, T57wx4, A67wx4, H67wx4, O67wx4, V67wx4, C77wx4;
wire J77wx4, Q77wx4, X77wx4, E87wx4, L87wx4, S87wx4, Z87wx4, G97wx4, N97wx4, U97wx4;
wire Ba7wx4, Ia7wx4, Pa7wx4, Wa7wx4, Db7wx4, Kb7wx4, Rb7wx4, Yb7wx4, Fc7wx4, Mc7wx4;
wire Tc7wx4, Ad7wx4, Hd7wx4, Od7wx4, Vd7wx4, Ce7wx4, Je7wx4, Qe7wx4, Xe7wx4, Ef7wx4;
wire Lf7wx4, Sf7wx4, Zf7wx4, Gg7wx4, Ng7wx4, Ug7wx4, Bh7wx4, Ih7wx4, Ph7wx4, Wh7wx4;
wire Di7wx4, Ki7wx4, Ri7wx4, Yi7wx4, Fj7wx4, Mj7wx4, Tj7wx4, Ak7wx4, Hk7wx4, Ok7wx4;
wire Vk7wx4, Cl7wx4, Jl7wx4, Ql7wx4, Xl7wx4, Em7wx4, Lm7wx4, Sm7wx4, Zm7wx4, Gn7wx4;
wire Nn7wx4, Un7wx4, Bo7wx4, Io7wx4, Po7wx4, Wo7wx4, Dp7wx4, Kp7wx4, Rp7wx4, Yp7wx4;
wire Fq7wx4, Mq7wx4, Tq7wx4, Ar7wx4, Hr7wx4, Or7wx4, Vr7wx4, Cs7wx4, Js7wx4, Qs7wx4;
wire Xs7wx4, Et7wx4, Lt7wx4, St7wx4, Zt7wx4, Gu7wx4, Nu7wx4, Uu7wx4, Bv7wx4, Iv7wx4;
wire Pv7wx4, Wv7wx4, Dw7wx4, Kw7wx4, Rw7wx4, Yw7wx4, Fx7wx4, Mx7wx4, Tx7wx4, Ay7wx4;
wire Hy7wx4, Oy7wx4, Vy7wx4, Cz7wx4, Jz7wx4, Qz7wx4, Xz7wx4, E08wx4, L08wx4, S08wx4;
wire Z08wx4, G18wx4, N18wx4, U18wx4, B28wx4, I28wx4, P28wx4, W28wx4, D38wx4, K38wx4;
wire R38wx4, Y38wx4, F48wx4, M48wx4, T48wx4, A58wx4, H58wx4, O58wx4, V58wx4, C68wx4;
wire J68wx4, Q68wx4, X68wx4, E78wx4, L78wx4, S78wx4, Z78wx4, G88wx4, N88wx4, U88wx4;
wire B98wx4, I98wx4, P98wx4, W98wx4, Da8wx4, Ka8wx4, Ra8wx4, Ya8wx4, Fb8wx4, Mb8wx4;
wire Tb8wx4, Ac8wx4, Hc8wx4, Oc8wx4, Vc8wx4, Cd8wx4, Jd8wx4, Qd8wx4, Xd8wx4, Ee8wx4;
wire Le8wx4, Se8wx4, Ze8wx4, Gf8wx4, Nf8wx4, Uf8wx4, Bg8wx4, Ig8wx4, Pg8wx4, Wg8wx4;
wire Dh8wx4, Kh8wx4, Rh8wx4, Yh8wx4, Fi8wx4, Mi8wx4, Ti8wx4, Aj8wx4, Hj8wx4, Oj8wx4;
wire Vj8wx4, Ck8wx4, Jk8wx4, Qk8wx4, Xk8wx4, El8wx4, Ll8wx4, Sl8wx4, Zl8wx4, Gm8wx4;
wire Nm8wx4, Um8wx4, Bn8wx4, In8wx4, Pn8wx4, Wn8wx4, Do8wx4, Ko8wx4, Ro8wx4, Yo8wx4;
wire Fp8wx4, Mp8wx4, Tp8wx4, Aq8wx4, Hq8wx4, Oq8wx4, Vq8wx4, Cr8wx4, Jr8wx4, Qr8wx4;
wire Xr8wx4, Es8wx4, Ls8wx4, Ss8wx4, Zs8wx4, Gt8wx4, Nt8wx4, Ut8wx4, Bu8wx4, Iu8wx4;
wire Pu8wx4, Wu8wx4, Dv8wx4, Kv8wx4, Rv8wx4, Yv8wx4, Fw8wx4, Mw8wx4, Tw8wx4, Ax8wx4;
wire Hx8wx4, Ox8wx4, Vx8wx4, Cy8wx4, Jy8wx4, Qy8wx4, Xy8wx4, Ez8wx4, Lz8wx4, Sz8wx4;
wire Zz8wx4, G09wx4, N09wx4, U09wx4, B19wx4, I19wx4, P19wx4, W19wx4, D29wx4, K29wx4;
wire R29wx4, Y29wx4, F39wx4, M39wx4, T39wx4, A49wx4, H49wx4, O49wx4, V49wx4, C59wx4;
wire J59wx4, Q59wx4, X59wx4, E69wx4, L69wx4, S69wx4, Z69wx4, G79wx4, N79wx4, U79wx4;
wire B89wx4, I89wx4, P89wx4, W89wx4, D99wx4, K99wx4, R99wx4, Y99wx4, Fa9wx4, Ma9wx4;
wire Ta9wx4, Ab9wx4, Hb9wx4, Ob9wx4, Vb9wx4, Cc9wx4, Jc9wx4, Qc9wx4, Xc9wx4, Ed9wx4;
wire Ld9wx4, Sd9wx4, Zd9wx4, Ge9wx4, Ne9wx4, Ue9wx4, Bf9wx4, If9wx4, Pf9wx4, Wf9wx4;
wire Dg9wx4, Kg9wx4, Rg9wx4, Yg9wx4, Fh9wx4, Mh9wx4, Th9wx4, Ai9wx4, Hi9wx4, Oi9wx4;
wire Vi9wx4, Cj9wx4, Jj9wx4, Qj9wx4, Xj9wx4, Ek9wx4, Lk9wx4, Sk9wx4, Zk9wx4, Gl9wx4;
wire Nl9wx4, Ul9wx4, Bm9wx4, Im9wx4, Pm9wx4, Wm9wx4, Dn9wx4, Kn9wx4, Rn9wx4, Yn9wx4;
wire Fo9wx4, Mo9wx4, To9wx4, Ap9wx4, Hp9wx4, Op9wx4, Vp9wx4, Cq9wx4, Jq9wx4, Qq9wx4;
wire Xq9wx4, Er9wx4, Lr9wx4, Sr9wx4, Zr9wx4, Gs9wx4, Ns9wx4, Us9wx4, Bt9wx4, It9wx4;
wire Pt9wx4, Wt9wx4, Du9wx4, Ku9wx4, Ru9wx4, Yu9wx4, Fv9wx4, Mv9wx4, Tv9wx4, Aw9wx4;
wire Hw9wx4, Ow9wx4, Vw9wx4, Cx9wx4, Jx9wx4, Qx9wx4, Xx9wx4, Ey9wx4, Ly9wx4, Sy9wx4;
wire Zy9wx4, Gz9wx4, Nz9wx4, Uz9wx4, B0awx4, I0awx4, P0awx4, W0awx4, D1awx4, K1awx4;
wire R1awx4, Y1awx4, F2awx4, M2awx4, T2awx4, A3awx4, H3awx4, O3awx4, V3awx4, C4awx4;
wire J4awx4, Q4awx4, X4awx4, E5awx4, L5awx4, S5awx4, Z5awx4, G6awx4, N6awx4, U6awx4;
wire B7awx4, I7awx4, P7awx4, W7awx4, D8awx4, K8awx4, R8awx4, Y8awx4, F9awx4, M9awx4;
wire T9awx4, Aaawx4, Haawx4, Oaawx4, Vaawx4, Cbawx4, Jbawx4, Qbawx4, Xbawx4, Ecawx4;
wire Lcawx4, Scawx4, Zcawx4, Gdawx4, Ndawx4, Udawx4, Beawx4, Ieawx4, Peawx4, Weawx4;
wire Dfawx4, Kfawx4, Rfawx4, Yfawx4, Fgawx4, Mgawx4, Tgawx4, Ahawx4, Hhawx4, Ohawx4;
wire Vhawx4, Ciawx4, Jiawx4, Qiawx4, Xiawx4, Ejawx4, Ljawx4, Sjawx4, Zjawx4, Gkawx4;
wire Nkawx4, Ukawx4, Blawx4, Ilawx4, Plawx4, Wlawx4, Dmawx4, Kmawx4, Rmawx4, Ymawx4;
wire Fnawx4, Mnawx4, Tnawx4, Aoawx4, Hoawx4, Ooawx4, Voawx4, Cpawx4, Jpawx4, Qpawx4;
wire Xpawx4, Eqawx4, Lqawx4, Sqawx4, Zqawx4, Grawx4, Nrawx4, Urawx4, Bsawx4, Isawx4;
wire Psawx4, Wsawx4, Dtawx4, Ktawx4, Rtawx4, Ytawx4, Fuawx4, Muawx4, Tuawx4, Avawx4;
wire Hvawx4, Ovawx4, Vvawx4, Cwawx4, Jwawx4, Qwawx4, Xwawx4, Exawx4, Lxawx4, Sxawx4;
wire Zxawx4, Gyawx4, Nyawx4, Uyawx4, Bzawx4, Izawx4, Pzawx4, Wzawx4, D0bwx4, K0bwx4;
wire R0bwx4, Y0bwx4, F1bwx4, M1bwx4, T1bwx4, A2bwx4, H2bwx4, O2bwx4, V2bwx4, C3bwx4;
wire J3bwx4, Q3bwx4, X3bwx4, E4bwx4, L4bwx4, S4bwx4, Z4bwx4, G5bwx4, N5bwx4, U5bwx4;
wire B6bwx4, I6bwx4, P6bwx4, W6bwx4, D7bwx4, K7bwx4, R7bwx4, Y7bwx4, F8bwx4, M8bwx4;
wire T8bwx4, A9bwx4, H9bwx4, O9bwx4, V9bwx4, Cabwx4, Jabwx4, Qabwx4, Xabwx4, Ebbwx4;
wire Lbbwx4, Sbbwx4, Zbbwx4, Gcbwx4, Ncbwx4, Ucbwx4, Bdbwx4, Idbwx4, Pdbwx4, Wdbwx4;
wire Debwx4, Kebwx4, Rebwx4, Yebwx4, Ffbwx4, Mfbwx4, Tfbwx4, Agbwx4, Hgbwx4, Ogbwx4;
wire Vgbwx4, Chbwx4, Jhbwx4, Qhbwx4, Xhbwx4, Eibwx4, Libwx4, Sibwx4, Zibwx4, Gjbwx4;
wire Njbwx4, Ujbwx4, Bkbwx4, Ikbwx4, Pkbwx4, Wkbwx4, Dlbwx4, Klbwx4, Rlbwx4, Ylbwx4;
wire Fmbwx4, Mmbwx4, Tmbwx4, Anbwx4, Hnbwx4, Onbwx4, Vnbwx4, Cobwx4, Jobwx4, Qobwx4;
wire Xobwx4, Epbwx4, Lpbwx4, Spbwx4, Zpbwx4, Gqbwx4, Nqbwx4, Uqbwx4, Brbwx4, Irbwx4;
wire Prbwx4, Wrbwx4, Dsbwx4, Ksbwx4, Rsbwx4, Ysbwx4, Ftbwx4, Mtbwx4, Ttbwx4, Aubwx4;
wire Hubwx4, Oubwx4, Vubwx4, Cvbwx4, Jvbwx4, Qvbwx4, Xvbwx4, Ewbwx4, Lwbwx4, Swbwx4;
wire Zwbwx4, Gxbwx4, Nxbwx4, Uxbwx4, Bybwx4, Iybwx4, Pybwx4, Wybwx4, Dzbwx4, Kzbwx4;
wire Rzbwx4, Yzbwx4, F0cwx4, M0cwx4, T0cwx4, A1cwx4, H1cwx4, O1cwx4, V1cwx4, C2cwx4;
wire J2cwx4, Q2cwx4, X2cwx4, E3cwx4, L3cwx4, S3cwx4, Z3cwx4, G4cwx4, N4cwx4, U4cwx4;
wire B5cwx4, I5cwx4, P5cwx4, W5cwx4, D6cwx4, K6cwx4, R6cwx4, Y6cwx4, F7cwx4, M7cwx4;
wire T7cwx4, A8cwx4, H8cwx4, O8cwx4, V8cwx4, C9cwx4, J9cwx4, Q9cwx4, X9cwx4, Eacwx4;
wire Lacwx4, Sacwx4, Zacwx4, Gbcwx4, Nbcwx4, Ubcwx4, Bccwx4, Iccwx4, Pccwx4, Wccwx4;
wire Ddcwx4, Kdcwx4, Rdcwx4, Ydcwx4, Fecwx4, Mecwx4, Tecwx4, Afcwx4, Hfcwx4, Ofcwx4;
wire Vfcwx4, Cgcwx4, Jgcwx4, Qgcwx4, Xgcwx4, Ehcwx4, Lhcwx4, Shcwx4, Zhcwx4, Gicwx4;
wire Nicwx4, Uicwx4, Bjcwx4, Ijcwx4, Pjcwx4, Wjcwx4, Dkcwx4, Kkcwx4, Rkcwx4, Ykcwx4;
wire Flcwx4, Mlcwx4, Tlcwx4, Amcwx4, Hmcwx4, Omcwx4, Vmcwx4, Cncwx4, Jncwx4, Qncwx4;
wire Xncwx4, Eocwx4, Locwx4, Socwx4, Zocwx4, Gpcwx4, Npcwx4, Upcwx4, Bqcwx4, Iqcwx4;
wire Pqcwx4, Wqcwx4, Drcwx4, Krcwx4, Rrcwx4, Yrcwx4, Fscwx4, Mscwx4, Tscwx4, Atcwx4;
wire Htcwx4, Otcwx4, Vtcwx4, Cucwx4, Jucwx4, Qucwx4, Xucwx4, Evcwx4, Lvcwx4, Svcwx4;
wire Zvcwx4, Gwcwx4, Nwcwx4, Uwcwx4, Bxcwx4, Ixcwx4, Pxcwx4, Wxcwx4, Dycwx4, Kycwx4;
wire Rycwx4, Yycwx4, Fzcwx4, Mzcwx4, Tzcwx4, A0dwx4, H0dwx4, O0dwx4, V0dwx4, C1dwx4;
wire J1dwx4, Q1dwx4, X1dwx4, E2dwx4, L2dwx4, S2dwx4, Z2dwx4, G3dwx4, N3dwx4, U3dwx4;
wire B4dwx4, I4dwx4, P4dwx4, W4dwx4, D5dwx4, K5dwx4, R5dwx4, Y5dwx4, F6dwx4, M6dwx4;
wire T6dwx4, A7dwx4, H7dwx4, O7dwx4, V7dwx4, C8dwx4, J8dwx4, Q8dwx4, X8dwx4, E9dwx4;
wire L9dwx4, S9dwx4, Z9dwx4, Gadwx4, Nadwx4, Uadwx4, Bbdwx4, Ibdwx4, Pbdwx4, Wbdwx4;
wire Dcdwx4, Kcdwx4, Rcdwx4, Ycdwx4, Fddwx4, Mddwx4, Tddwx4, Aedwx4, Hedwx4, Oedwx4;
wire Vedwx4, Cfdwx4, Jfdwx4, Qfdwx4, Xfdwx4, Egdwx4, Lgdwx4, Sgdwx4, Zgdwx4, Ghdwx4;
wire Nhdwx4, Uhdwx4, Bidwx4, Iidwx4, Pidwx4, Widwx4, Djdwx4, Kjdwx4, Rjdwx4, Yjdwx4;
wire Fkdwx4, Mkdwx4, Tkdwx4, Aldwx4, Hldwx4, Oldwx4, Vldwx4, Cmdwx4, Jmdwx4, Qmdwx4;
wire Xmdwx4, Endwx4, Lndwx4, Sndwx4, Zndwx4, Godwx4, Nodwx4, Uodwx4, Bpdwx4, Ipdwx4;
wire Ppdwx4, Wpdwx4, Dqdwx4, Kqdwx4, Rqdwx4, Yqdwx4, Frdwx4, Mrdwx4, Trdwx4, Asdwx4;
wire Hsdwx4, Osdwx4, Vsdwx4, Ctdwx4, Jtdwx4, Qtdwx4, Xtdwx4, Eudwx4, Ludwx4, Sudwx4;
wire Zudwx4, Gvdwx4, Nvdwx4, Uvdwx4, Bwdwx4, Iwdwx4, Pwdwx4, Wwdwx4, Dxdwx4, Kxdwx4;
wire Rxdwx4, Yxdwx4, Fydwx4, Mydwx4, Tydwx4, Azdwx4, Hzdwx4, Ozdwx4, Vzdwx4, C0ewx4;
wire J0ewx4, Q0ewx4, X0ewx4, E1ewx4, L1ewx4, S1ewx4, Z1ewx4, G2ewx4, N2ewx4, U2ewx4;
wire B3ewx4, I3ewx4, P3ewx4, W3ewx4, D4ewx4, K4ewx4, R4ewx4, Y4ewx4, F5ewx4, M5ewx4;
wire T5ewx4, A6ewx4, H6ewx4, O6ewx4, V6ewx4, C7ewx4, J7ewx4, Q7ewx4, X7ewx4, E8ewx4;
wire L8ewx4, S8ewx4, Z8ewx4, G9ewx4, N9ewx4, U9ewx4, Baewx4, Iaewx4, Paewx4, Waewx4;
wire Dbewx4, Kbewx4, Rbewx4, Ybewx4, Fcewx4, Mcewx4, Tcewx4, Adewx4, Hdewx4, Odewx4;
wire Vdewx4, Ceewx4, Jeewx4, Qeewx4, Xeewx4, Efewx4, Lfewx4, Sfewx4, Zfewx4, Ggewx4;
wire Ngewx4, Ugewx4, Bhewx4, Ihewx4, Phewx4, Whewx4, Diewx4, Kiewx4, Riewx4, Yiewx4;
wire Fjewx4, Mjewx4, Tjewx4, Akewx4, Hkewx4, Okewx4, Vkewx4, Clewx4, Jlewx4, Qlewx4;
wire Xlewx4, Emewx4, Lmewx4, Smewx4, Zmewx4, Gnewx4, Nnewx4, Unewx4, Boewx4, Ioewx4;
wire Poewx4, Woewx4, Dpewx4, Kpewx4, Rpewx4, Ypewx4, Fqewx4, Mqewx4, Tqewx4, Arewx4;
wire Hrewx4, Orewx4, Vrewx4, Csewx4, Jsewx4, Qsewx4, Xsewx4, Etewx4, Ltewx4, Stewx4;
wire Ztewx4, Guewx4, Nuewx4, Uuewx4, Bvewx4, Ivewx4, Pvewx4, Wvewx4, Dwewx4, Kwewx4;
wire Rwewx4, Ywewx4, Fxewx4, Mxewx4, Txewx4, Ayewx4, Hyewx4, Oyewx4, Vyewx4, Czewx4;
wire Jzewx4, Qzewx4, Xzewx4, E0fwx4, L0fwx4, S0fwx4, Z0fwx4, G1fwx4, N1fwx4, U1fwx4;
wire B2fwx4, I2fwx4, P2fwx4, W2fwx4, D3fwx4, K3fwx4, R3fwx4, Y3fwx4, F4fwx4, M4fwx4;
wire T4fwx4, A5fwx4, H5fwx4, O5fwx4, V5fwx4, C6fwx4, J6fwx4, Q6fwx4, X6fwx4, E7fwx4;
wire L7fwx4, S7fwx4, Z7fwx4, G8fwx4, N8fwx4, U8fwx4, B9fwx4, I9fwx4, P9fwx4, W9fwx4;
wire Dafwx4, Kafwx4, Rafwx4, Yafwx4, Fbfwx4, Mbfwx4, Tbfwx4, Acfwx4, Hcfwx4, Ocfwx4;
wire Vcfwx4, Cdfwx4, Jdfwx4, Qdfwx4, Xdfwx4, Eefwx4, Lefwx4, Sefwx4, Zefwx4, Gffwx4;
wire Nffwx4, Uffwx4, Bgfwx4, Igfwx4, Pgfwx4, Wgfwx4, Dhfwx4, Khfwx4, Rhfwx4, Yhfwx4;
wire Fifwx4, Mifwx4, Tifwx4, Ajfwx4, Hjfwx4, Ojfwx4, Vjfwx4, Ckfwx4, Jkfwx4, Qkfwx4;
wire Xkfwx4, Elfwx4, Llfwx4, Slfwx4, Zlfwx4, Gmfwx4, Nmfwx4, Umfwx4, Bnfwx4, Infwx4;
wire Pnfwx4, Wnfwx4, Dofwx4, Kofwx4, Rofwx4, Yofwx4, Fpfwx4, Mpfwx4, Tpfwx4, Aqfwx4;
wire Hqfwx4, Oqfwx4, Vqfwx4, Crfwx4, Jrfwx4, Qrfwx4, Xrfwx4, Esfwx4, Lsfwx4, Ssfwx4;
wire Zsfwx4, Gtfwx4, Ntfwx4, Utfwx4, Bufwx4, Iufwx4, Pufwx4, Wufwx4, Dvfwx4, Kvfwx4;
wire Rvfwx4, Yvfwx4, Fwfwx4, Mwfwx4, Twfwx4, Axfwx4, Hxfwx4, Oxfwx4, Vxfwx4, Cyfwx4;
wire Jyfwx4, Qyfwx4, Xyfwx4, Ezfwx4, Lzfwx4, Szfwx4, Zzfwx4, G0gwx4, N0gwx4, U0gwx4;
wire B1gwx4, I1gwx4, P1gwx4, W1gwx4, D2gwx4, K2gwx4, R2gwx4, Y2gwx4, F3gwx4, M3gwx4;
wire T3gwx4, A4gwx4, H4gwx4, O4gwx4, V4gwx4, C5gwx4, J5gwx4, Q5gwx4, X5gwx4, E6gwx4;
wire L6gwx4, S6gwx4, Z6gwx4, G7gwx4, N7gwx4, U7gwx4, B8gwx4, I8gwx4, P8gwx4, W8gwx4;
wire D9gwx4, K9gwx4, R9gwx4, Y9gwx4, Fagwx4, Magwx4, Tagwx4, Abgwx4, Hbgwx4, Obgwx4;
wire Vbgwx4, Ccgwx4, Jcgwx4, Qcgwx4, Xcgwx4, Edgwx4, Ldgwx4, Sdgwx4, Zdgwx4, Gegwx4;
wire Negwx4, Uegwx4, Bfgwx4, Ifgwx4, Pfgwx4, Wfgwx4, Dggwx4, Kggwx4, Rggwx4, Yggwx4;
wire Fhgwx4, Mhgwx4, Thgwx4, Aigwx4, Higwx4, Oigwx4, Vigwx4, Cjgwx4, Jjgwx4, Qjgwx4;
wire Xjgwx4, Ekgwx4, Lkgwx4, Skgwx4, Zkgwx4, Glgwx4, Nlgwx4, Ulgwx4, Bmgwx4, Imgwx4;
wire Pmgwx4, Wmgwx4, Dngwx4, Kngwx4, Rngwx4, Yngwx4, Fogwx4, Mogwx4, Togwx4, Apgwx4;
wire Hpgwx4, Opgwx4, Vpgwx4, Cqgwx4, Jqgwx4, Qqgwx4, Xqgwx4, Ergwx4, Lrgwx4, Srgwx4;
wire Zrgwx4, Gsgwx4, Nsgwx4, Usgwx4, Btgwx4, Itgwx4, Ptgwx4, Wtgwx4, Dugwx4, Kugwx4;
wire Rugwx4, Yugwx4, Fvgwx4, Mvgwx4, Tvgwx4, Awgwx4, Hwgwx4, Owgwx4, Vwgwx4, Cxgwx4;
wire Jxgwx4, Qxgwx4, Xxgwx4, Eygwx4, Lygwx4, Sygwx4, Zygwx4, Gzgwx4, Nzgwx4, Uzgwx4;
wire B0hwx4, I0hwx4, P0hwx4, W0hwx4, D1hwx4, K1hwx4, R1hwx4, Y1hwx4, F2hwx4, M2hwx4;
wire T2hwx4, A3hwx4, H3hwx4, O3hwx4, V3hwx4, C4hwx4, J4hwx4, Q4hwx4, X4hwx4, E5hwx4;
wire L5hwx4, S5hwx4, Z5hwx4, G6hwx4, N6hwx4, U6hwx4, B7hwx4, I7hwx4, P7hwx4, W7hwx4;
wire D8hwx4, K8hwx4, R8hwx4, Y8hwx4, F9hwx4, M9hwx4, T9hwx4, Aahwx4, Hahwx4, Oahwx4;
wire Vahwx4, Cbhwx4, Jbhwx4, Qbhwx4, Xbhwx4, Echwx4, Lchwx4, Schwx4, Zchwx4, Gdhwx4;
wire Ndhwx4, Udhwx4, Behwx4, Iehwx4, Pehwx4, Wehwx4, Dfhwx4, Kfhwx4, Rfhwx4, Yfhwx4;
wire Fghwx4, Mghwx4, Tghwx4, Ahhwx4, Hhhwx4, Ohhwx4, Vhhwx4, Cihwx4, Jihwx4, Qihwx4;
wire Xihwx4, Ejhwx4, Ljhwx4, Sjhwx4, Zjhwx4, Gkhwx4, Nkhwx4, Ukhwx4, Blhwx4, Ilhwx4;
wire Plhwx4, Wlhwx4, Dmhwx4, Kmhwx4, Rmhwx4, Ymhwx4, Fnhwx4, Mnhwx4, Tnhwx4, Aohwx4;
wire Hohwx4, Oohwx4, Vohwx4, Cphwx4, Jphwx4, Qphwx4, Xphwx4, Eqhwx4, Lqhwx4, Sqhwx4;
wire Zqhwx4, Grhwx4, Nrhwx4, Urhwx4, Bshwx4, Ishwx4, Pshwx4, Wshwx4, Dthwx4, Kthwx4;
wire Rthwx4, Ythwx4, Fuhwx4, Muhwx4, Tuhwx4, Avhwx4, Hvhwx4, Ovhwx4, Vvhwx4, Cwhwx4;
wire Jwhwx4, Qwhwx4, Xwhwx4, Exhwx4, Lxhwx4, Sxhwx4, Zxhwx4, Gyhwx4, Nyhwx4, Uyhwx4;
wire Bzhwx4, Izhwx4, Pzhwx4, Wzhwx4, D0iwx4, K0iwx4, R0iwx4, Y0iwx4, F1iwx4, M1iwx4;
wire T1iwx4, A2iwx4, H2iwx4, O2iwx4, V2iwx4, C3iwx4, J3iwx4, Q3iwx4, X3iwx4, E4iwx4;
wire L4iwx4, S4iwx4, Z4iwx4, G5iwx4, N5iwx4, U5iwx4, B6iwx4, I6iwx4, P6iwx4, W6iwx4;
wire D7iwx4, K7iwx4, R7iwx4, Y7iwx4, F8iwx4, M8iwx4, T8iwx4, A9iwx4, H9iwx4, O9iwx4;
wire V9iwx4, Caiwx4, Jaiwx4, Qaiwx4, Xaiwx4, Ebiwx4, Lbiwx4, Sbiwx4, Zbiwx4, Gciwx4;
wire Nciwx4, Uciwx4, Bdiwx4, Idiwx4, Pdiwx4, Wdiwx4, Deiwx4, Keiwx4, Reiwx4, Yeiwx4;
wire Ffiwx4, Mfiwx4, Tfiwx4, Agiwx4, Hgiwx4, Ogiwx4, Vgiwx4, Chiwx4, Jhiwx4, Qhiwx4;
wire Xhiwx4, Eiiwx4, Liiwx4, Siiwx4, Ziiwx4, Gjiwx4, Njiwx4, Ujiwx4, Bkiwx4, Ikiwx4;
wire Pkiwx4, Wkiwx4, Dliwx4, Kliwx4, Rliwx4, Yliwx4, Fmiwx4, Mmiwx4, Tmiwx4, Aniwx4;
wire Hniwx4, Oniwx4, Vniwx4, Coiwx4, Joiwx4, Qoiwx4, Xoiwx4, Epiwx4, Lpiwx4, Spiwx4;
wire Zpiwx4, Gqiwx4, Nqiwx4, Uqiwx4, Briwx4, Iriwx4, Priwx4, Wriwx4, Dsiwx4, Ksiwx4;
wire Rsiwx4, Ysiwx4, Ftiwx4, Mtiwx4, Ttiwx4, Auiwx4, Huiwx4, Ouiwx4, Vuiwx4, Cviwx4;
wire Jviwx4, Qviwx4, Xviwx4, Ewiwx4, Lwiwx4, Swiwx4, Zwiwx4, Gxiwx4, Nxiwx4, Uxiwx4;
wire Byiwx4, Iyiwx4, Pyiwx4, Wyiwx4, Dziwx4, Kziwx4, Rziwx4, Yziwx4, F0jwx4, M0jwx4;
wire T0jwx4, A1jwx4, H1jwx4, O1jwx4, V1jwx4, C2jwx4, J2jwx4, Q2jwx4, X2jwx4, E3jwx4;
wire L3jwx4, S3jwx4, Z3jwx4, G4jwx4, N4jwx4, U4jwx4, B5jwx4, I5jwx4, P5jwx4, W5jwx4;
wire D6jwx4, K6jwx4, R6jwx4, Y6jwx4, F7jwx4, M7jwx4, T7jwx4, A8jwx4, H8jwx4, O8jwx4;
wire V8jwx4, C9jwx4, J9jwx4, Q9jwx4, X9jwx4, Eajwx4, Lajwx4, Sajwx4, Zajwx4, Gbjwx4;
wire Nbjwx4, Ubjwx4, Bcjwx4, Icjwx4, Pcjwx4, Wcjwx4, Ddjwx4, Kdjwx4, Rdjwx4, Ydjwx4;
wire Fejwx4, Mejwx4, Tejwx4, Afjwx4, Hfjwx4, Ofjwx4, Vfjwx4, Cgjwx4, Jgjwx4, Qgjwx4;
wire Xgjwx4, Ehjwx4, Lhjwx4, Shjwx4, Zhjwx4, Gijwx4, Nijwx4, Uijwx4, Bjjwx4, Ijjwx4;
wire Pjjwx4, Wjjwx4, Dkjwx4, Kkjwx4, Rkjwx4, Ykjwx4, Fljwx4, Mljwx4, Tljwx4, Amjwx4;
wire Hmjwx4, Omjwx4, Vmjwx4, Cnjwx4, Jnjwx4, Qnjwx4, Xnjwx4, Eojwx4, Lojwx4, Sojwx4;
wire Zojwx4, Gpjwx4, Npjwx4, Upjwx4, Bqjwx4, Iqjwx4, Pqjwx4, Wqjwx4, Drjwx4, Krjwx4;
wire Rrjwx4, Yrjwx4, Fsjwx4, Msjwx4, Tsjwx4, Atjwx4, Htjwx4, Otjwx4, Vtjwx4, Cujwx4;
wire Jujwx4, Qujwx4, Xujwx4, Evjwx4, Lvjwx4, Svjwx4, Zvjwx4, Gwjwx4, Nwjwx4, Uwjwx4;
wire Bxjwx4, Ixjwx4, Pxjwx4, Wxjwx4, Dyjwx4, Kyjwx4, Ryjwx4, Yyjwx4, Fzjwx4, Mzjwx4;
wire Tzjwx4, A0kwx4, H0kwx4, O0kwx4, V0kwx4, C1kwx4, J1kwx4, Q1kwx4, X1kwx4, E2kwx4;
wire L2kwx4, S2kwx4, Z2kwx4, G3kwx4, N3kwx4, U3kwx4, B4kwx4, I4kwx4, P4kwx4, W4kwx4;
wire D5kwx4, K5kwx4, R5kwx4, Y5kwx4, F6kwx4, M6kwx4, T6kwx4, A7kwx4, H7kwx4, O7kwx4;
wire V7kwx4, C8kwx4, J8kwx4, Q8kwx4, X8kwx4, E9kwx4, L9kwx4, S9kwx4, Z9kwx4, Gakwx4;
wire Nakwx4, Uakwx4, Bbkwx4, Ibkwx4, Pbkwx4, Wbkwx4, Dckwx4, Kckwx4, Rckwx4, Yckwx4;
wire Fdkwx4, Mdkwx4, Tdkwx4, Aekwx4, Hekwx4, Oekwx4, Vekwx4, Cfkwx4, Jfkwx4, Qfkwx4;
wire Xfkwx4, Egkwx4, Lgkwx4, Sgkwx4, Zgkwx4, Ghkwx4, Nhkwx4, Uhkwx4, Bikwx4, Iikwx4;
wire Pikwx4, Wikwx4, Djkwx4, Kjkwx4, Rjkwx4, Yjkwx4, Fkkwx4, Mkkwx4, Tkkwx4, Alkwx4;
wire Hlkwx4, Olkwx4, Vlkwx4, Cmkwx4, Jmkwx4, Qmkwx4, Xmkwx4, Enkwx4, Lnkwx4, Snkwx4;
wire Znkwx4, Gokwx4, Nokwx4, Uokwx4, Bpkwx4, Ipkwx4, Ppkwx4, Wpkwx4, Dqkwx4, Kqkwx4;
wire Rqkwx4, Yqkwx4, Frkwx4, Mrkwx4, Trkwx4, Askwx4, Hskwx4, Oskwx4, Vskwx4, Ctkwx4;
wire Jtkwx4, Qtkwx4, Xtkwx4, Eukwx4, Lukwx4, Sukwx4, Zukwx4, Gvkwx4, Nvkwx4, Uvkwx4;
wire Bwkwx4, Iwkwx4, Pwkwx4, Wwkwx4, Dxkwx4, Kxkwx4, Rxkwx4, Yxkwx4, Fykwx4, Mykwx4;
wire Tykwx4, Azkwx4, Hzkwx4, Ozkwx4, Vzkwx4, C0lwx4, J0lwx4, Q0lwx4, X0lwx4, E1lwx4;
wire L1lwx4, S1lwx4, Z1lwx4, G2lwx4, N2lwx4, U2lwx4, B3lwx4, I3lwx4, P3lwx4, W3lwx4;
wire D4lwx4, K4lwx4, R4lwx4, Y4lwx4, F5lwx4, M5lwx4, T5lwx4, A6lwx4, H6lwx4, O6lwx4;
wire V6lwx4, C7lwx4, J7lwx4, Q7lwx4, X7lwx4, E8lwx4, L8lwx4, S8lwx4, Z8lwx4, G9lwx4;
wire N9lwx4, U9lwx4, Balwx4, Ialwx4, Palwx4, Walwx4, Dblwx4, Kblwx4, Rblwx4, Yblwx4;
wire Fclwx4, Mclwx4, Tclwx4, Adlwx4, Hdlwx4, Odlwx4, Vdlwx4, Celwx4, Jelwx4, Qelwx4;
wire Xelwx4, Eflwx4, Lflwx4, Sflwx4, Zflwx4, Gglwx4, Nglwx4, Uglwx4, Bhlwx4, Ihlwx4;
wire Phlwx4, Whlwx4, Dilwx4, Kilwx4, Rilwx4, Yilwx4, Fjlwx4, Mjlwx4, Tjlwx4, Aklwx4;
wire Hklwx4, Oklwx4, Vklwx4, Cllwx4, Jllwx4, Qllwx4, Xllwx4, Emlwx4, Lmlwx4, Smlwx4;
wire Zmlwx4, Gnlwx4, Nnlwx4, Unlwx4, Bolwx4, Iolwx4, Polwx4, Wolwx4, Dplwx4, Kplwx4;
wire Rplwx4, Yplwx4, Fqlwx4, Mqlwx4, Tqlwx4, Arlwx4, Hrlwx4, Orlwx4, Vrlwx4, Cslwx4;
wire Jslwx4, Qslwx4, Xslwx4, Etlwx4, Ltlwx4, Stlwx4, Ztlwx4, Gulwx4, Nulwx4, Uulwx4;
wire Bvlwx4, Ivlwx4, Pvlwx4, Wvlwx4, Dwlwx4, Kwlwx4, Rwlwx4, Ywlwx4, Fxlwx4, Mxlwx4;
wire Txlwx4, Aylwx4, Hylwx4, Oylwx4, Vylwx4, Czlwx4, Jzlwx4, Qzlwx4, Xzlwx4, E0mwx4;
wire L0mwx4, S0mwx4, Z0mwx4, G1mwx4, N1mwx4, U1mwx4, B2mwx4, I2mwx4, P2mwx4, W2mwx4;
wire D3mwx4, K3mwx4, R3mwx4, Y3mwx4, F4mwx4, M4mwx4, T4mwx4, A5mwx4, H5mwx4, O5mwx4;
wire V5mwx4, C6mwx4, J6mwx4, Q6mwx4, X6mwx4, E7mwx4, L7mwx4, S7mwx4, Z7mwx4, G8mwx4;
wire N8mwx4, U8mwx4, B9mwx4, I9mwx4, P9mwx4, W9mwx4, Damwx4, Kamwx4, Ramwx4, Yamwx4;
wire Fbmwx4, Mbmwx4, Tbmwx4, Acmwx4, Hcmwx4, Ocmwx4, Vcmwx4, Cdmwx4, Jdmwx4, Qdmwx4;
wire Xdmwx4, Eemwx4, Lemwx4, Semwx4, Zemwx4, Gfmwx4, Nfmwx4, Ufmwx4, Bgmwx4, Igmwx4;
wire Pgmwx4, Wgmwx4, Dhmwx4, Khmwx4, Rhmwx4, Yhmwx4, Fimwx4, Mimwx4, Timwx4, Ajmwx4;
wire Hjmwx4, Ojmwx4, Vjmwx4, Ckmwx4, Jkmwx4, Qkmwx4, Xkmwx4, Elmwx4, Llmwx4, Slmwx4;
wire Zlmwx4, Gmmwx4, Nmmwx4, Ummwx4, Bnmwx4, Inmwx4, Pnmwx4, Wnmwx4, Domwx4, Komwx4;
wire Romwx4, Yomwx4, Fpmwx4, Mpmwx4, Tpmwx4, Aqmwx4, Hqmwx4, Oqmwx4, Vqmwx4, Crmwx4;
wire Jrmwx4, Qrmwx4, Xrmwx4, Esmwx4, Lsmwx4, Ssmwx4, Zsmwx4, Gtmwx4, Ntmwx4, Utmwx4;
wire Bumwx4, Iumwx4, Pumwx4, Wumwx4, Dvmwx4, Kvmwx4, Rvmwx4, Yvmwx4, Fwmwx4, Mwmwx4;
wire Twmwx4, Axmwx4, Hxmwx4, Oxmwx4, Vxmwx4, Cymwx4, Jymwx4, Qymwx4, Xymwx4, Ezmwx4;
wire Lzmwx4, Szmwx4, Zzmwx4, G0nwx4, N0nwx4, U0nwx4, B1nwx4, I1nwx4, P1nwx4, W1nwx4;
wire D2nwx4, K2nwx4, R2nwx4, Y2nwx4, F3nwx4, M3nwx4, T3nwx4, A4nwx4, H4nwx4, O4nwx4;
wire V4nwx4, C5nwx4, J5nwx4, Q5nwx4, X5nwx4, E6nwx4, L6nwx4, S6nwx4, Z6nwx4, G7nwx4;
wire N7nwx4, U7nwx4, B8nwx4, I8nwx4, P8nwx4, W8nwx4, D9nwx4, K9nwx4, R9nwx4, Y9nwx4;
wire Fanwx4, Manwx4, Tanwx4, Abnwx4, Hbnwx4, Obnwx4, Vbnwx4, Ccnwx4, Jcnwx4, Qcnwx4;
wire Xcnwx4, Ednwx4, Ldnwx4, Sdnwx4, Zdnwx4, Genwx4, Nenwx4, Uenwx4, Bfnwx4, Ifnwx4;
wire Pfnwx4, Wfnwx4, Dgnwx4, Kgnwx4, Rgnwx4, Ygnwx4, Fhnwx4, Mhnwx4, Thnwx4, Ainwx4;
wire Hinwx4, Oinwx4, Vinwx4, Cjnwx4, Jjnwx4, Qjnwx4, Xjnwx4, Eknwx4, Lknwx4, Sknwx4;
wire Zknwx4, Glnwx4, Nlnwx4, Ulnwx4, Bmnwx4, Imnwx4, Pmnwx4, Wmnwx4, Dnnwx4, Knnwx4;
wire Rnnwx4, Ynnwx4, Fonwx4, Monwx4, Tonwx4, Apnwx4, Hpnwx4, Opnwx4, Vpnwx4, Cqnwx4;
wire Jqnwx4, Qqnwx4, Xqnwx4, Ernwx4, Lrnwx4, Srnwx4, Zrnwx4, Gsnwx4, Nsnwx4, Usnwx4;
wire Btnwx4, Itnwx4, Ptnwx4, Wtnwx4, Dunwx4, Kunwx4, Runwx4, Yunwx4, Fvnwx4, Mvnwx4;
wire Tvnwx4, Awnwx4, Hwnwx4, Ownwx4, Vwnwx4, Cxnwx4, Jxnwx4, Qxnwx4, Xxnwx4, Eynwx4;
wire Lynwx4, Synwx4, Zynwx4, Gznwx4, Nznwx4, Uznwx4, B0owx4, I0owx4, P0owx4, W0owx4;
wire D1owx4, K1owx4, R1owx4, Y1owx4, F2owx4, M2owx4, T2owx4, A3owx4, H3owx4, O3owx4;
wire V3owx4, C4owx4, J4owx4, Q4owx4, X4owx4, E5owx4, L5owx4, S5owx4, Z5owx4, G6owx4;
wire N6owx4, U6owx4, B7owx4, I7owx4, P7owx4, W7owx4, D8owx4, K8owx4, R8owx4, Y8owx4;
wire F9owx4, M9owx4, T9owx4, Aaowx4, Haowx4, Oaowx4, Vaowx4, Cbowx4, Jbowx4, Qbowx4;
wire Xbowx4, Ecowx4, Lcowx4, Scowx4, Zcowx4, Gdowx4, Ndowx4, Udowx4, Beowx4, Ieowx4;
wire Peowx4, Weowx4, Dfowx4, Kfowx4, Rfowx4, Yfowx4, Fgowx4, Mgowx4, Tgowx4, Ahowx4;
wire Hhowx4, Ohowx4, Vhowx4, Ciowx4, Jiowx4, Qiowx4, Xiowx4, Ejowx4, Ljowx4, Sjowx4;
wire Zjowx4, Gkowx4, Nkowx4, Ukowx4, Blowx4, Ilowx4, Plowx4, Wlowx4, Dmowx4, Kmowx4;
wire Rmowx4, Ymowx4, Fnowx4, Mnowx4, Tnowx4, Aoowx4, Hoowx4, Ooowx4, Voowx4, Cpowx4;
wire Jpowx4, Qpowx4, Xpowx4, Eqowx4, Lqowx4, Sqowx4, Zqowx4, Growx4, Nrowx4, Urowx4;
wire Bsowx4, Isowx4, Psowx4, Wsowx4, Dtowx4, Ktowx4, Rtowx4, Ytowx4, Fuowx4, Muowx4;
wire Tuowx4, Avowx4, Hvowx4, Ovowx4, Vvowx4, Cwowx4, Jwowx4, Qwowx4, Xwowx4, Exowx4;
wire Lxowx4, Sxowx4, Zxowx4, Gyowx4, Nyowx4, Uyowx4, Bzowx4, Izowx4, Pzowx4, Wzowx4;
wire D0pwx4, K0pwx4, R0pwx4, Y0pwx4, F1pwx4, M1pwx4, T1pwx4, A2pwx4, H2pwx4, O2pwx4;
wire V2pwx4, C3pwx4, J3pwx4, Q3pwx4, X3pwx4, E4pwx4, L4pwx4, S4pwx4, Z4pwx4, G5pwx4;
wire N5pwx4, U5pwx4, B6pwx4, I6pwx4, P6pwx4, W6pwx4, D7pwx4, K7pwx4, R7pwx4, Y7pwx4;
wire F8pwx4, M8pwx4, T8pwx4, A9pwx4, H9pwx4, O9pwx4, V9pwx4, Capwx4, Japwx4, Qapwx4;
wire Xapwx4, Ebpwx4, Lbpwx4, Sbpwx4, Zbpwx4, Gcpwx4, Ncpwx4, Ucpwx4, Bdpwx4, Idpwx4;
wire Pdpwx4, Wdpwx4, Depwx4, Kepwx4, Repwx4, Yepwx4, Ffpwx4, Mfpwx4, Tfpwx4, Agpwx4;
wire Hgpwx4, Ogpwx4, Vgpwx4, Chpwx4, Jhpwx4, Qhpwx4, Xhpwx4, Eipwx4, Lipwx4, Sipwx4;
wire Zipwx4, Gjpwx4, Njpwx4, Ujpwx4, Bkpwx4, Ikpwx4, Pkpwx4, Wkpwx4, Dlpwx4, Klpwx4;
wire Rlpwx4, Ylpwx4, Fmpwx4, Mmpwx4, Tmpwx4, Anpwx4, Hnpwx4, Onpwx4, Vnpwx4, Copwx4;
wire Jopwx4, Qopwx4, Xopwx4, Eppwx4, Lppwx4, Sppwx4, Zppwx4, Gqpwx4, Nqpwx4, Uqpwx4;
wire Brpwx4, Irpwx4, Prpwx4, Wrpwx4, Dspwx4, Kspwx4, Rspwx4, Yspwx4, Ftpwx4, Mtpwx4;
wire Ttpwx4, Aupwx4, Hupwx4, Oupwx4, Vupwx4, Cvpwx4, Jvpwx4, Qvpwx4, Xvpwx4, Ewpwx4;
wire Lwpwx4, Swpwx4, Zwpwx4, Gxpwx4, Nxpwx4, Uxpwx4, Bypwx4, Iypwx4, Pypwx4, Wypwx4;
wire Dzpwx4, Kzpwx4, Rzpwx4, Yzpwx4, F0qwx4, M0qwx4, T0qwx4, A1qwx4, H1qwx4, O1qwx4;
wire V1qwx4, C2qwx4, J2qwx4, Q2qwx4, X2qwx4, E3qwx4, L3qwx4, S3qwx4, Z3qwx4, G4qwx4;
wire N4qwx4, U4qwx4, B5qwx4, I5qwx4, P5qwx4, W5qwx4, D6qwx4, K6qwx4, R6qwx4, Y6qwx4;
wire F7qwx4, M7qwx4, T7qwx4, A8qwx4, H8qwx4, O8qwx4, V8qwx4, C9qwx4, J9qwx4, Q9qwx4;
wire X9qwx4, Eaqwx4, Laqwx4, Saqwx4, Zaqwx4, Gbqwx4, Nbqwx4, Ubqwx4, Bcqwx4, Icqwx4;
wire Pcqwx4, Wcqwx4, Ddqwx4, Kdqwx4, Rdqwx4, Ydqwx4, Feqwx4, Meqwx4, Teqwx4, Afqwx4;
wire Hfqwx4, Ofqwx4, Vfqwx4, Cgqwx4, Jgqwx4, Qgqwx4, Xgqwx4, Ehqwx4, Lhqwx4, Shqwx4;
wire Zhqwx4, Giqwx4, Niqwx4, Uiqwx4, Bjqwx4, Ijqwx4, Pjqwx4, Wjqwx4, Dkqwx4, Kkqwx4;
wire Rkqwx4, Ykqwx4, Flqwx4, Mlqwx4, Tlqwx4, Amqwx4, Hmqwx4, Omqwx4, Vmqwx4, Cnqwx4;
wire Jnqwx4, Qnqwx4, Xnqwx4, Eoqwx4, Loqwx4, Soqwx4, Zoqwx4, Gpqwx4, Npqwx4, Upqwx4;
wire Bqqwx4, Iqqwx4, Pqqwx4, Wqqwx4, Drqwx4, Krqwx4, Rrqwx4, Yrqwx4, Fsqwx4, Msqwx4;
wire Tsqwx4, Atqwx4, Htqwx4, Otqwx4, Vtqwx4, Cuqwx4, Juqwx4, Quqwx4, Xuqwx4, Evqwx4;
wire Lvqwx4, Svqwx4, Zvqwx4, Gwqwx4, Nwqwx4, Uwqwx4, Bxqwx4, Ixqwx4, Pxqwx4, Wxqwx4;
wire Dyqwx4, Kyqwx4, Ryqwx4, Yyqwx4, Fzqwx4, Mzqwx4, Tzqwx4, A0rwx4, H0rwx4, O0rwx4;
wire V0rwx4, C1rwx4, J1rwx4, Q1rwx4, X1rwx4, E2rwx4, L2rwx4, S2rwx4, Z2rwx4, G3rwx4;
wire N3rwx4, U3rwx4, B4rwx4, I4rwx4, P4rwx4, W4rwx4, D5rwx4, K5rwx4, R5rwx4, Y5rwx4;
wire F6rwx4, M6rwx4, T6rwx4, A7rwx4, H7rwx4, O7rwx4, V7rwx4, C8rwx4, J8rwx4, Q8rwx4;
wire X8rwx4, E9rwx4, L9rwx4, S9rwx4, Z9rwx4, Garwx4, Narwx4, Uarwx4, Bbrwx4, Ibrwx4;
wire Pbrwx4, Wbrwx4, Dcrwx4, Kcrwx4, Rcrwx4, Ycrwx4, Fdrwx4, Mdrwx4, Tdrwx4, Aerwx4;
wire Herwx4, Oerwx4, Verwx4, Cfrwx4, Jfrwx4, Qfrwx4, Xfrwx4, Egrwx4, Lgrwx4, Sgrwx4;
wire Zgrwx4, Ghrwx4, Nhrwx4, Uhrwx4, Birwx4, Iirwx4, Pirwx4, Wirwx4, Djrwx4, Kjrwx4;
wire Rjrwx4, Yjrwx4, Fkrwx4, Mkrwx4, Tkrwx4, Alrwx4, Hlrwx4, Olrwx4, Vlrwx4, Cmrwx4;
wire Jmrwx4, Qmrwx4, Xmrwx4, Enrwx4, Lnrwx4, Snrwx4, Znrwx4, Gorwx4, Norwx4, Uorwx4;
wire Bprwx4, Iprwx4, Pprwx4, Wprwx4, Dqrwx4, Kqrwx4, Rqrwx4, Yqrwx4, Frrwx4, Mrrwx4;
wire Trrwx4, Asrwx4, Hsrwx4, Osrwx4, Vsrwx4, Ctrwx4, Jtrwx4, Qtrwx4, Xtrwx4, Eurwx4;
wire Lurwx4, Surwx4, Zurwx4, Gvrwx4, Nvrwx4, Uvrwx4, Bwrwx4, Iwrwx4, Pwrwx4, Wwrwx4;
wire Dxrwx4, Kxrwx4, Rxrwx4, Yxrwx4, Fyrwx4, Myrwx4, Tyrwx4, Azrwx4, Hzrwx4, Ozrwx4;
wire Vzrwx4, C0swx4, J0swx4, Q0swx4, X0swx4, E1swx4, L1swx4, S1swx4, Z1swx4, G2swx4;
wire N2swx4, U2swx4, B3swx4, I3swx4, P3swx4, W3swx4, D4swx4, K4swx4, R4swx4, Y4swx4;
wire F5swx4, M5swx4, T5swx4, A6swx4, H6swx4, O6swx4, V6swx4, C7swx4, J7swx4, Q7swx4;
wire X7swx4, E8swx4, L8swx4, S8swx4, Z8swx4, G9swx4, N9swx4, U9swx4, Baswx4, Iaswx4;
wire Paswx4, Waswx4, Dbswx4, Kbswx4, Rbswx4, Ybswx4, Fcswx4, Mcswx4, Tcswx4, Adswx4;
wire Hdswx4, Odswx4, Vdswx4, Ceswx4, Jeswx4, Qeswx4, Xeswx4, Efswx4, Lfswx4, Sfswx4;
wire Zfswx4, Ggswx4, Ngswx4, Ugswx4, Bhswx4, Ihswx4, Phswx4, Whswx4, Diswx4, Kiswx4;
wire Riswx4, Yiswx4, Fjswx4, Mjswx4, Tjswx4, Akswx4, Hkswx4, Okswx4, Vkswx4, Clswx4;
wire Jlswx4, Qlswx4, Xlswx4, Emswx4, Lmswx4, Smswx4, Zmswx4, Gnswx4, Nnswx4, Unswx4;
wire Boswx4, Ioswx4, Poswx4, Woswx4, Dpswx4, Kpswx4, Rpswx4, Ypswx4, Fqswx4, Mqswx4;
wire Tqswx4, Arswx4, Hrswx4, Orswx4, Vrswx4, Csswx4, Jsswx4, Qsswx4, Xsswx4, Etswx4;
wire Ltswx4, Stswx4, Ztswx4, Guswx4, Nuswx4, Uuswx4, Bvswx4, Ivswx4, Pvswx4, Wvswx4;
wire Dwswx4, Kwswx4, Rwswx4, Ywswx4, Fxswx4, Mxswx4, Txswx4, Ayswx4, Hyswx4, Oyswx4;
wire Vyswx4, Czswx4, Jzswx4, Qzswx4, Xzswx4, E0twx4, L0twx4, S0twx4, Z0twx4, G1twx4;
wire N1twx4, U1twx4, B2twx4, I2twx4, P2twx4, W2twx4, D3twx4, K3twx4, R3twx4, Y3twx4;
wire F4twx4, M4twx4, T4twx4, A5twx4, H5twx4, O5twx4, V5twx4, C6twx4, J6twx4, Q6twx4;
wire X6twx4, E7twx4, L7twx4, S7twx4, Z7twx4, G8twx4, N8twx4, U8twx4, B9twx4, I9twx4;
wire P9twx4, W9twx4, Datwx4, Katwx4, Ratwx4, Yatwx4, Fbtwx4, Mbtwx4, Tbtwx4, Actwx4;
wire Hctwx4, Octwx4, Vctwx4, Cdtwx4, Jdtwx4, Qdtwx4, Xdtwx4, Eetwx4, Letwx4, Setwx4;
wire Zetwx4, Gftwx4, Nftwx4, Uftwx4, Bgtwx4, Igtwx4, Pgtwx4, Wgtwx4, Dhtwx4, Khtwx4;
wire Rhtwx4, Yhtwx4, Fitwx4, Mitwx4, Titwx4, Ajtwx4, Hjtwx4, Ojtwx4, Vjtwx4, Cktwx4;
wire Jktwx4, Qktwx4, Xktwx4, Eltwx4, Lltwx4, Sltwx4, Zltwx4, Gmtwx4, Nmtwx4, Umtwx4;
wire Bntwx4, Intwx4, Pntwx4, Wntwx4, Dotwx4, Kotwx4, Rotwx4, Yotwx4, Fptwx4, Mptwx4;
wire Tptwx4, Aqtwx4, Hqtwx4, Oqtwx4, Vqtwx4, Crtwx4, Jrtwx4, Qrtwx4, Xrtwx4, Estwx4;
wire Lstwx4, Sstwx4, Zstwx4, Gttwx4, Nttwx4, Uttwx4, Butwx4, Iutwx4, Putwx4, Wutwx4;
wire Dvtwx4, Kvtwx4, Rvtwx4, Yvtwx4, Fwtwx4, Mwtwx4, Twtwx4, Axtwx4, Hxtwx4, Oxtwx4;
wire Vxtwx4, Cytwx4, Jytwx4, Qytwx4, Xytwx4, Eztwx4, Lztwx4, Sztwx4, Zztwx4, G0uwx4;
wire N0uwx4, U0uwx4, B1uwx4, I1uwx4, P1uwx4, W1uwx4, D2uwx4, K2uwx4, R2uwx4, Y2uwx4;
wire F3uwx4, M3uwx4, T3uwx4, A4uwx4, H4uwx4, O4uwx4, V4uwx4, C5uwx4, J5uwx4, Q5uwx4;
wire X5uwx4, E6uwx4, L6uwx4, S6uwx4, Z6uwx4, G7uwx4, N7uwx4, U7uwx4, B8uwx4, I8uwx4;
wire P8uwx4, W8uwx4, D9uwx4, K9uwx4, R9uwx4, Y9uwx4, Fauwx4, Mauwx4, Tauwx4, Abuwx4;
wire Hbuwx4, Obuwx4, Vbuwx4, Ccuwx4, Jcuwx4, Qcuwx4, Xcuwx4, Eduwx4, Lduwx4, Sduwx4;
wire Zduwx4, Geuwx4, Neuwx4, Ueuwx4, Bfuwx4, Ifuwx4, Pfuwx4, Wfuwx4, Dguwx4, Kguwx4;
wire Rguwx4, Yguwx4, Fhuwx4, Mhuwx4, Thuwx4, Aiuwx4, Hiuwx4, Oiuwx4, Viuwx4, Cjuwx4;
wire Jjuwx4, Qjuwx4, Xjuwx4, Ekuwx4, Lkuwx4, Skuwx4, Zkuwx4, Gluwx4, Nluwx4, Uluwx4;
wire Bmuwx4, Imuwx4, Pmuwx4, Wmuwx4, Dnuwx4, Knuwx4, Rnuwx4, Ynuwx4, Fouwx4, Mouwx4;
wire Touwx4, Apuwx4, Hpuwx4, Opuwx4, Vpuwx4, Cquwx4, Jquwx4, Qquwx4, Xquwx4, Eruwx4;
wire Lruwx4, Sruwx4, Zruwx4, Gsuwx4, Nsuwx4, Usuwx4, Btuwx4, Ituwx4, Ptuwx4, Wtuwx4;
wire Duuwx4, Kuuwx4, Ruuwx4, Yuuwx4, Fvuwx4, Mvuwx4, Tvuwx4, Awuwx4, Hwuwx4, Owuwx4;
wire Vwuwx4, Cxuwx4, Jxuwx4, Qxuwx4, Xxuwx4, Eyuwx4, Lyuwx4, Syuwx4, Zyuwx4, Gzuwx4;
wire Nzuwx4, Uzuwx4, B0vwx4, I0vwx4, P0vwx4, W0vwx4, D1vwx4, K1vwx4, R1vwx4, Y1vwx4;
wire F2vwx4, M2vwx4, T2vwx4, A3vwx4, H3vwx4, O3vwx4, V3vwx4, C4vwx4, J4vwx4, Q4vwx4;
wire X4vwx4, E5vwx4, L5vwx4, S5vwx4, Z5vwx4, G6vwx4, N6vwx4, U6vwx4, B7vwx4, I7vwx4;
wire P7vwx4, W7vwx4, D8vwx4, K8vwx4, R8vwx4, Y8vwx4, F9vwx4, M9vwx4, T9vwx4, Aavwx4;
wire Havwx4, Oavwx4, Vavwx4, Cbvwx4, Jbvwx4, Qbvwx4, Xbvwx4, Ecvwx4, Lcvwx4, Scvwx4;
wire Zcvwx4, Gdvwx4, Ndvwx4, Udvwx4, Bevwx4, Ievwx4, Pevwx4, Wevwx4, Dfvwx4, Kfvwx4;
wire Rfvwx4, Yfvwx4, Fgvwx4, Mgvwx4, Tgvwx4, Ahvwx4, Hhvwx4, Ohvwx4, Vhvwx4, Civwx4;
wire Jivwx4, Qivwx4, Xivwx4, Ejvwx4, Ljvwx4, Sjvwx4, Zjvwx4, Gkvwx4, Nkvwx4, Ukvwx4;
wire Blvwx4, Ilvwx4, Plvwx4, Wlvwx4, Dmvwx4, Kmvwx4, Rmvwx4, Ymvwx4, Fnvwx4, Mnvwx4;
wire Tnvwx4, Aovwx4, Hovwx4, Oovwx4, Vovwx4, Cpvwx4, Jpvwx4, Qpvwx4, Xpvwx4, Eqvwx4;
wire Lqvwx4, Sqvwx4, Zqvwx4, Grvwx4, Nrvwx4, Urvwx4, Bsvwx4, Isvwx4, Psvwx4, Wsvwx4;
wire Dtvwx4, Ktvwx4, Rtvwx4, Ytvwx4, Fuvwx4, Muvwx4, Tuvwx4, Avvwx4, Hvvwx4, Ovvwx4;
wire Vvvwx4, Cwvwx4, Jwvwx4, Qwvwx4, Xwvwx4, Exvwx4, Lxvwx4, Sxvwx4, Zxvwx4, Gyvwx4;
wire Nyvwx4, Uyvwx4, Bzvwx4, Izvwx4, Pzvwx4, Wzvwx4, D0wwx4, K0wwx4, R0wwx4, Y0wwx4;
wire F1wwx4, M1wwx4, T1wwx4, A2wwx4, H2wwx4, O2wwx4, V2wwx4, C3wwx4, J3wwx4, Q3wwx4;
wire X3wwx4, E4wwx4, L4wwx4, S4wwx4, Z4wwx4, G5wwx4, N5wwx4, U5wwx4, B6wwx4, I6wwx4;
wire P6wwx4, W6wwx4, D7wwx4, K7wwx4, R7wwx4, Y7wwx4, F8wwx4, M8wwx4, T8wwx4, A9wwx4;
wire H9wwx4, O9wwx4, V9wwx4, Cawwx4, Jawwx4, Qawwx4, Xawwx4, Ebwwx4, Lbwwx4, Sbwwx4;
wire Zbwwx4, Gcwwx4, Ncwwx4, Ucwwx4, Bdwwx4, Idwwx4, Pdwwx4, Wdwwx4, Dewwx4, Kewwx4;
wire Rewwx4, Yewwx4, Ffwwx4, Mfwwx4, Tfwwx4, Agwwx4, Hgwwx4, Ogwwx4, Vgwwx4, Chwwx4;
wire Jhwwx4, Qhwwx4, Xhwwx4, Eiwwx4, Liwwx4, Siwwx4, Ziwwx4, Gjwwx4, Njwwx4, Ujwwx4;
wire Bkwwx4, Ikwwx4, Pkwwx4, Wkwwx4, Dlwwx4, Klwwx4, Rlwwx4, Ylwwx4, Fmwwx4, Mmwwx4;
wire Tmwwx4, Anwwx4, Hnwwx4, Onwwx4, Vnwwx4, Cowwx4, Jowwx4, Qowwx4, Xowwx4, Epwwx4;
wire Lpwwx4, Spwwx4, Zpwwx4, Gqwwx4, Nqwwx4, Uqwwx4, Brwwx4, Irwwx4, Prwwx4, Wrwwx4;
wire Dswwx4, Kswwx4, Rswwx4, Yswwx4, Ftwwx4, Mtwwx4, Ttwwx4, Auwwx4, Huwwx4, Ouwwx4;
wire Vuwwx4, Cvwwx4, Jvwwx4, Qvwwx4, Xvwwx4, Ewwwx4, Lwwwx4, Swwwx4, Zwwwx4, Gxwwx4;
wire Nxwwx4, Uxwwx4, Bywwx4, Iywwx4, Pywwx4, Wywwx4, Dzwwx4, Kzwwx4, Rzwwx4, Yzwwx4;
wire F0xwx4, M0xwx4, T0xwx4, A1xwx4, H1xwx4, O1xwx4, V1xwx4, C2xwx4, J2xwx4, Q2xwx4;
wire X2xwx4, E3xwx4, L3xwx4, S3xwx4, Z3xwx4, G4xwx4, N4xwx4, U4xwx4, B5xwx4, I5xwx4;
wire P5xwx4, W5xwx4, D6xwx4, K6xwx4, R6xwx4, Y6xwx4, F7xwx4, M7xwx4, T7xwx4, A8xwx4;
wire H8xwx4, O8xwx4, V8xwx4, C9xwx4, J9xwx4, Q9xwx4, X9xwx4, Eaxwx4, Laxwx4, Saxwx4;
wire Zaxwx4, Gbxwx4, Nbxwx4, Ubxwx4, Bcxwx4, Icxwx4, Pcxwx4, Wcxwx4, Ddxwx4, Kdxwx4;
wire Rdxwx4, Ydxwx4, Fexwx4, Mexwx4, Texwx4, Afxwx4, Hfxwx4, Ofxwx4, Vfxwx4, Cgxwx4;
wire Jgxwx4, Qgxwx4, Xgxwx4, Ehxwx4, Lhxwx4, Shxwx4, Zhxwx4, Gixwx4, Nixwx4, Uixwx4;
wire Bjxwx4, Ijxwx4, Pjxwx4, Wjxwx4, Dkxwx4, Kkxwx4, Rkxwx4, Ykxwx4, Flxwx4, Mlxwx4;
wire Tlxwx4, Amxwx4, Hmxwx4, Omxwx4, Vmxwx4, Cnxwx4, Jnxwx4, Qnxwx4, Xnxwx4, Eoxwx4;
wire Loxwx4, Soxwx4, Zoxwx4, Gpxwx4, Npxwx4, Upxwx4, Bqxwx4, Iqxwx4, Pqxwx4, Wqxwx4;
wire Drxwx4, Krxwx4, Rrxwx4, Yrxwx4, Fsxwx4, Msxwx4, Tsxwx4, Atxwx4, Htxwx4, Otxwx4;
wire Vtxwx4, Cuxwx4, Juxwx4, Quxwx4, Xuxwx4, Evxwx4, Lvxwx4, Svxwx4, Zvxwx4, Gwxwx4;
wire Nwxwx4, Uwxwx4, Bxxwx4, Ixxwx4, Pxxwx4, Wxxwx4, Dyxwx4, Kyxwx4, Ryxwx4, Yyxwx4;
wire Fzxwx4, Mzxwx4, Tzxwx4, A0ywx4, H0ywx4, O0ywx4, V0ywx4, C1ywx4, J1ywx4, Q1ywx4;
wire X1ywx4, E2ywx4, L2ywx4, S2ywx4, Z2ywx4, G3ywx4, N3ywx4, U3ywx4, B4ywx4, I4ywx4;
wire P4ywx4, W4ywx4, D5ywx4, K5ywx4, R5ywx4, Y5ywx4, F6ywx4, M6ywx4, T6ywx4, A7ywx4;
wire H7ywx4, O7ywx4, V7ywx4, C8ywx4, J8ywx4, Q8ywx4, X8ywx4, E9ywx4, L9ywx4, S9ywx4;
wire Z9ywx4, Gaywx4, Naywx4, Uaywx4, Bbywx4, Ibywx4, Pbywx4, Wbywx4, Dcywx4, Kcywx4;
wire Rcywx4, Ycywx4, Fdywx4, Mdywx4, Tdywx4, Aeywx4, Heywx4, Oeywx4, Veywx4, Cfywx4;
wire Jfywx4, Qfywx4, Xfywx4, Egywx4, Lgywx4, Sgywx4, Zgywx4, Ghywx4, Nhywx4, Uhywx4;
wire Biywx4, Iiywx4, Piywx4, Wiywx4, Djywx4, Kjywx4, Rjywx4, Yjywx4, Fkywx4, Mkywx4;
wire Tkywx4, Alywx4, Hlywx4, Olywx4, Vlywx4, Cmywx4, Jmywx4, Qmywx4, Xmywx4, Enywx4;
wire Lnywx4, Snywx4, Znywx4, Goywx4, Noywx4, Uoywx4, Bpywx4, Ipywx4, Ppywx4, Wpywx4;
wire Dqywx4, Kqywx4, Rqywx4, Yqywx4, Frywx4, Mrywx4, Trywx4, Asywx4, Hsywx4, Osywx4;
wire Vsywx4, Ctywx4, Jtywx4, Qtywx4, Xtywx4, Euywx4, Luywx4, Suywx4, Zuywx4, Gvywx4;
wire Nvywx4, Uvywx4, Bwywx4, Iwywx4, Pwywx4, Wwywx4, Dxywx4, Kxywx4, Rxywx4, Yxywx4;
wire Fyywx4, Myywx4, Tyywx4, Azywx4, Hzywx4, Ozywx4, Vzywx4, C0zwx4, J0zwx4, Q0zwx4;
wire X0zwx4, E1zwx4, L1zwx4, S1zwx4, Z1zwx4, G2zwx4, N2zwx4, U2zwx4, B3zwx4, I3zwx4;
wire P3zwx4, W3zwx4, D4zwx4, K4zwx4, R4zwx4, Y4zwx4, F5zwx4, M5zwx4, T5zwx4, A6zwx4;
wire H6zwx4, O6zwx4, V6zwx4, C7zwx4, J7zwx4, Q7zwx4, X7zwx4, E8zwx4, L8zwx4, S8zwx4;
wire Z8zwx4, G9zwx4, N9zwx4, U9zwx4, Bazwx4, Iazwx4, Pazwx4, Wazwx4, Dbzwx4, Kbzwx4;
wire Rbzwx4, Ybzwx4, Fczwx4, Mczwx4, Tczwx4, Adzwx4, Hdzwx4, Odzwx4, Vdzwx4, Cezwx4;
wire Jezwx4, Qezwx4, Xezwx4, Efzwx4, Lfzwx4, Sfzwx4, Zfzwx4, Ggzwx4, Ngzwx4, Ugzwx4;
wire Bhzwx4, Ihzwx4, Phzwx4, Whzwx4, Dizwx4, Kizwx4, Rizwx4, Yizwx4, Fjzwx4, Mjzwx4;
wire Tjzwx4, Akzwx4, Hkzwx4, Okzwx4, Vkzwx4, Clzwx4, Jlzwx4, Qlzwx4, Xlzwx4, Emzwx4;
wire Lmzwx4, Smzwx4, Zmzwx4, Gnzwx4, Nnzwx4, Unzwx4, Bozwx4, Iozwx4, Pozwx4, Wozwx4;
wire Dpzwx4, Kpzwx4, Rpzwx4, Ypzwx4, Fqzwx4, Mqzwx4, Tqzwx4, Arzwx4, Hrzwx4, Orzwx4;
wire Vrzwx4, Cszwx4, Jszwx4, Qszwx4, Xszwx4, Etzwx4, Ltzwx4, Stzwx4, Ztzwx4, Guzwx4;
wire Nuzwx4, Uuzwx4, Bvzwx4, Ivzwx4, Pvzwx4, Wvzwx4, Dwzwx4, Kwzwx4, Rwzwx4, Ywzwx4;
wire Fxzwx4, Mxzwx4, Txzwx4, Ayzwx4, Hyzwx4, Oyzwx4, Vyzwx4, Czzwx4, Jzzwx4, Qzzwx4;
wire Xzzwx4, E00xx4, L00xx4, S00xx4, Z00xx4, G10xx4, N10xx4, U10xx4, B20xx4, I20xx4;
wire P20xx4, W20xx4, D30xx4, K30xx4, R30xx4, Y30xx4, F40xx4, M40xx4, T40xx4, A50xx4;
wire H50xx4, O50xx4, V50xx4, C60xx4, J60xx4, Q60xx4, X60xx4, E70xx4, L70xx4, S70xx4;
wire Z70xx4, G80xx4, N80xx4, U80xx4, B90xx4, I90xx4, P90xx4, W90xx4, Da0xx4, Ka0xx4;
wire Ra0xx4, Ya0xx4, Fb0xx4, Mb0xx4, Tb0xx4, Ac0xx4, Hc0xx4, Oc0xx4, Vc0xx4, Cd0xx4;
wire Jd0xx4, Qd0xx4, Xd0xx4, Ee0xx4, Le0xx4, Se0xx4, Ze0xx4, Gf0xx4, Nf0xx4, Uf0xx4;
wire Bg0xx4, Ig0xx4, Pg0xx4, Wg0xx4, Dh0xx4, Kh0xx4, Rh0xx4, Yh0xx4, Fi0xx4, Mi0xx4;
wire Ti0xx4, Aj0xx4, Hj0xx4, Oj0xx4, Vj0xx4, Ck0xx4, Jk0xx4, Qk0xx4, Xk0xx4, El0xx4;
wire Ll0xx4, Sl0xx4, Zl0xx4, Gm0xx4, Nm0xx4, Um0xx4, Bn0xx4, In0xx4, Pn0xx4, Wn0xx4;
wire Do0xx4, Ko0xx4, Ro0xx4, Yo0xx4, Fp0xx4, Mp0xx4, Tp0xx4, Aq0xx4, Hq0xx4, Oq0xx4;
wire Vq0xx4, Cr0xx4, Jr0xx4, Qr0xx4, Xr0xx4, Es0xx4, Ls0xx4, Ss0xx4, Zs0xx4, Gt0xx4;
wire Nt0xx4, Ut0xx4, Bu0xx4, Iu0xx4, Pu0xx4, Wu0xx4, Dv0xx4, Kv0xx4, Rv0xx4, Yv0xx4;
wire Fw0xx4, Mw0xx4, Tw0xx4, Ax0xx4, Hx0xx4, Ox0xx4, Vx0xx4, Cy0xx4, Jy0xx4, Qy0xx4;
wire Xy0xx4, Ez0xx4, Lz0xx4, Sz0xx4, Zz0xx4, G01xx4, N01xx4, U01xx4, B11xx4, I11xx4;
wire P11xx4, W11xx4, D21xx4, K21xx4, R21xx4, Y21xx4, F31xx4, M31xx4, T31xx4, A41xx4;
wire H41xx4, O41xx4, V41xx4, C51xx4, J51xx4, Q51xx4, X51xx4, E61xx4, L61xx4, S61xx4;
wire Z61xx4, G71xx4, N71xx4, U71xx4, B81xx4, I81xx4, P81xx4, W81xx4, D91xx4, K91xx4;
wire R91xx4, Y91xx4, Fa1xx4, Ma1xx4, Ta1xx4, Ab1xx4, Hb1xx4, Ob1xx4, Vb1xx4, Cc1xx4;
wire Jc1xx4, Qc1xx4, Xc1xx4, Ed1xx4, Ld1xx4, Sd1xx4, Zd1xx4, Ge1xx4, Ne1xx4, Ue1xx4;
wire Bf1xx4, If1xx4, Pf1xx4, Wf1xx4, Dg1xx4, Kg1xx4, Rg1xx4, Yg1xx4, Fh1xx4, Mh1xx4;
wire Th1xx4, Ai1xx4, Hi1xx4, Oi1xx4, Vi1xx4, Cj1xx4, Jj1xx4, Qj1xx4, Xj1xx4, Ek1xx4;
wire Lk1xx4, Sk1xx4, Zk1xx4, Gl1xx4, Nl1xx4, Ul1xx4, Bm1xx4, Im1xx4, Pm1xx4, Wm1xx4;
wire Dn1xx4, Kn1xx4, Rn1xx4, Yn1xx4, Fo1xx4, Mo1xx4, To1xx4, Ap1xx4, Hp1xx4, Op1xx4;
wire Vp1xx4, Cq1xx4, Jq1xx4, Qq1xx4, Xq1xx4, Er1xx4, Lr1xx4, Sr1xx4, Zr1xx4, Gs1xx4;
wire Ns1xx4, Us1xx4, Bt1xx4, It1xx4, Pt1xx4, Wt1xx4, Du1xx4, Ku1xx4, Ru1xx4, Yu1xx4;
wire Fv1xx4, Mv1xx4, Tv1xx4, Aw1xx4, Hw1xx4, Ow1xx4, Vw1xx4, Cx1xx4, Jx1xx4, Qx1xx4;
wire Xx1xx4, Ey1xx4, Ly1xx4, Sy1xx4, Zy1xx4, Gz1xx4, Nz1xx4, Uz1xx4, B02xx4, I02xx4;
wire P02xx4, W02xx4, D12xx4, K12xx4, R12xx4, Y12xx4, F22xx4, M22xx4, T22xx4, A32xx4;
wire H32xx4, O32xx4, V32xx4, C42xx4, J42xx4, Q42xx4, X42xx4, E52xx4, L52xx4, S52xx4;
wire Z52xx4, G62xx4, N62xx4, U62xx4, B72xx4, I72xx4, P72xx4, W72xx4, D82xx4, K82xx4;
wire R82xx4, Y82xx4, F92xx4, M92xx4, T92xx4, Aa2xx4, Ha2xx4, Oa2xx4, Va2xx4, Cb2xx4;
wire Jb2xx4, Qb2xx4, Xb2xx4, Ec2xx4, Lc2xx4, Sc2xx4, Zc2xx4, Gd2xx4, Nd2xx4, Ud2xx4;
wire Be2xx4, Ie2xx4, Pe2xx4, We2xx4, Df2xx4, Kf2xx4, Rf2xx4, Yf2xx4, Fg2xx4, Mg2xx4;
wire Tg2xx4, Ah2xx4, Hh2xx4, Oh2xx4, Vh2xx4, Ci2xx4, Ji2xx4, Qi2xx4, Xi2xx4, Ej2xx4;
wire Lj2xx4, Sj2xx4, Zj2xx4, Gk2xx4, Nk2xx4, Uk2xx4, Bl2xx4, Il2xx4, Pl2xx4, Wl2xx4;
wire Dm2xx4, Km2xx4, Rm2xx4, Ym2xx4, Fn2xx4, Mn2xx4, Tn2xx4, Ao2xx4, Ho2xx4, Oo2xx4;
wire Vo2xx4, Cp2xx4, Jp2xx4, Qp2xx4, Xp2xx4, Eq2xx4, Lq2xx4, Sq2xx4, Zq2xx4, Gr2xx4;
wire Nr2xx4, Ur2xx4, Bs2xx4, Is2xx4, Ps2xx4, Ws2xx4, Dt2xx4, Kt2xx4, Rt2xx4, Yt2xx4;
wire Fu2xx4, Mu2xx4, Tu2xx4, Av2xx4, Hv2xx4, Ov2xx4, Vv2xx4, Cw2xx4, Jw2xx4, Qw2xx4;
wire Xw2xx4, Ex2xx4, Lx2xx4, Sx2xx4, Zx2xx4, Gy2xx4, Ny2xx4, Uy2xx4, Bz2xx4, Iz2xx4;
wire Pz2xx4, Wz2xx4, D03xx4, K03xx4, R03xx4, Y03xx4, F13xx4, M13xx4, T13xx4, A23xx4;
wire H23xx4, O23xx4, V23xx4, C33xx4, J33xx4, Q33xx4, X33xx4, E43xx4, L43xx4, S43xx4;
wire Z43xx4, G53xx4, N53xx4, U53xx4, B63xx4, I63xx4, P63xx4, W63xx4, D73xx4, K73xx4;
wire R73xx4, Y73xx4, F83xx4, M83xx4, T83xx4, A93xx4, H93xx4, O93xx4, V93xx4, Ca3xx4;
wire Ja3xx4, Qa3xx4, Xa3xx4, Eb3xx4, Lb3xx4, Sb3xx4, Zb3xx4, Gc3xx4, Nc3xx4, Uc3xx4;
wire Bd3xx4, Id3xx4, Pd3xx4, Wd3xx4, De3xx4, Ke3xx4, Re3xx4, Ye3xx4, Ff3xx4, Mf3xx4;
wire Tf3xx4, Ag3xx4, Hg3xx4, Og3xx4, Vg3xx4, Ch3xx4, Jh3xx4, Qh3xx4, Xh3xx4, Ei3xx4;
wire Li3xx4, Si3xx4, Zi3xx4, Gj3xx4, Nj3xx4, Uj3xx4, Bk3xx4, Ik3xx4, Pk3xx4, Wk3xx4;
wire Dl3xx4, Kl3xx4, Rl3xx4, Yl3xx4, Fm3xx4, Mm3xx4, Tm3xx4, An3xx4, Hn3xx4, On3xx4;
wire Vn3xx4, Co3xx4, Jo3xx4, Qo3xx4, Xo3xx4, Ep3xx4, Lp3xx4, Sp3xx4, Zp3xx4, Gq3xx4;
wire Nq3xx4, Uq3xx4, Br3xx4, Ir3xx4, Pr3xx4, Wr3xx4, Ds3xx4, Ks3xx4, Rs3xx4, Ys3xx4;
wire Ft3xx4, Mt3xx4, Tt3xx4, Au3xx4, Hu3xx4, Ou3xx4, Vu3xx4, Cv3xx4, Jv3xx4, Qv3xx4;
wire Xv3xx4, Ew3xx4, Lw3xx4, Sw3xx4, Zw3xx4, Gx3xx4, Nx3xx4, Ux3xx4, By3xx4, Iy3xx4;
wire Py3xx4, Wy3xx4, Dz3xx4, Kz3xx4, Rz3xx4, Yz3xx4, F04xx4, M04xx4, T04xx4, A14xx4;
wire H14xx4, O14xx4, V14xx4, C24xx4, J24xx4, Q24xx4, X24xx4, E34xx4, L34xx4, S34xx4;
wire Z34xx4, G44xx4, N44xx4, U44xx4, B54xx4, I54xx4, P54xx4, W54xx4, D64xx4, K64xx4;
wire R64xx4, Y64xx4, F74xx4, M74xx4, T74xx4, A84xx4, H84xx4, O84xx4, V84xx4, C94xx4;
wire J94xx4, Q94xx4, X94xx4, Ea4xx4, La4xx4, Sa4xx4, Za4xx4, Gb4xx4, Nb4xx4, Ub4xx4;
wire Bc4xx4, Ic4xx4, Pc4xx4, Wc4xx4, Dd4xx4, Kd4xx4, Rd4xx4, Yd4xx4, Fe4xx4, Me4xx4;
wire Te4xx4, Af4xx4, Hf4xx4, Of4xx4, Vf4xx4, Cg4xx4, Jg4xx4, Qg4xx4, Xg4xx4, Eh4xx4;
wire Lh4xx4, Sh4xx4, Zh4xx4, Gi4xx4, Ni4xx4, Ui4xx4, Bj4xx4, Ij4xx4, Pj4xx4, Wj4xx4;
wire Dk4xx4, Kk4xx4, Rk4xx4, Yk4xx4, Fl4xx4, Ml4xx4, Tl4xx4, Am4xx4, Hm4xx4, Om4xx4;
wire Vm4xx4, Cn4xx4, Jn4xx4, Qn4xx4, Xn4xx4, Eo4xx4, Lo4xx4, So4xx4, Zo4xx4, Gp4xx4;
wire Np4xx4, Up4xx4, Bq4xx4, Iq4xx4, Pq4xx4, Wq4xx4, Dr4xx4, Kr4xx4, Rr4xx4, Yr4xx4;
wire Fs4xx4, Ms4xx4, Ts4xx4, At4xx4, Ht4xx4, Ot4xx4, Vt4xx4, Cu4xx4, Ju4xx4, Qu4xx4;
wire Xu4xx4, Ev4xx4, Lv4xx4, Sv4xx4, Zv4xx4, Gw4xx4, Nw4xx4, Uw4xx4, Bx4xx4, Ix4xx4;
wire Px4xx4, Wx4xx4, Dy4xx4, Ky4xx4, Ry4xx4, Yy4xx4, Fz4xx4, Mz4xx4, Tz4xx4, A05xx4;
wire H05xx4, O05xx4, V05xx4, C15xx4, J15xx4, Q15xx4, X15xx4, E25xx4, L25xx4, S25xx4;
wire Z25xx4, G35xx4, N35xx4, U35xx4, B45xx4, I45xx4, P45xx4, W45xx4, D55xx4, K55xx4;
wire R55xx4, Y55xx4, F65xx4, M65xx4, T65xx4, A75xx4, H75xx4, O75xx4, V75xx4, C85xx4;
wire J85xx4, Q85xx4, X85xx4, E95xx4, L95xx4, S95xx4, Z95xx4, Ga5xx4, Na5xx4, Ua5xx4;
wire Bb5xx4, Ib5xx4, Pb5xx4, Wb5xx4, Dc5xx4, Kc5xx4, Rc5xx4, Yc5xx4, Fd5xx4, Md5xx4;
wire Td5xx4, Ae5xx4, He5xx4, Oe5xx4, Ve5xx4, Cf5xx4, Jf5xx4, Qf5xx4, Xf5xx4, Eg5xx4;
wire Lg5xx4, Sg5xx4, Zg5xx4, Gh5xx4, Nh5xx4, Uh5xx4, Bi5xx4, Ii5xx4, Pi5xx4, Wi5xx4;
wire Dj5xx4, Kj5xx4, Rj5xx4, Yj5xx4, Fk5xx4, Mk5xx4, Tk5xx4, Al5xx4, Hl5xx4, Ol5xx4;
wire Vl5xx4, Cm5xx4, Jm5xx4, Qm5xx4, Xm5xx4, En5xx4, Ln5xx4, Sn5xx4, Zn5xx4, Go5xx4;
wire No5xx4, Uo5xx4, Bp5xx4, Ip5xx4, Pp5xx4, Wp5xx4, Dq5xx4, Kq5xx4, Rq5xx4, Yq5xx4;
wire Fr5xx4, Mr5xx4, Tr5xx4, As5xx4, Hs5xx4, Os5xx4, Vs5xx4, Ct5xx4, Jt5xx4, Qt5xx4;
wire Xt5xx4, Eu5xx4, Lu5xx4, Su5xx4, Zu5xx4, Gv5xx4, Nv5xx4, Uv5xx4, Bw5xx4, Iw5xx4;
wire Pw5xx4, Ww5xx4, Dx5xx4, Ol22z4, Vl22z4, Cm22z4, Jm22z4, Qm22z4, Xm22z4, En22z4;
wire Ln22z4, Sn22z4, Zn22z4, Go22z4, No22z4, Uo22z4, Bp22z4, Ip22z4, Pp22z4, Wp22z4;
wire Dq22z4, Kq22z4, Rq22z4, Yq22z4, Fr22z4, Mr22z4, Tr22z4, As22z4, Hs22z4, Os22z4;
wire Vs22z4, Ct22z4, Jt22z4, Qt22z4, Xt22z4, Eu22z4, Lu22z4, Su22z4, Zu22z4, Gv22z4;
wire Nv22z4, Uv22z4, Bw22z4, Iw22z4, Pw22z4, Ww22z4, Dx22z4, Kx22z4, Rx22z4, Yx22z4;
wire Fy22z4, My22z4, Ty22z4, Az22z4, Hz22z4, Oz22z4, Vz22z4, C032z4, J032z4, Q032z4;
wire X032z4, E132z4, L132z4, S132z4, Z132z4, G232z4, N232z4, U232z4, B332z4, I332z4;
wire P332z4, W332z4, D432z4, K432z4, R432z4, Y432z4, F532z4, M532z4, T532z4, A632z4;
wire H632z4, O632z4, V632z4, C732z4, J732z4, Q732z4, X732z4, E832z4, L832z4, S832z4;
wire Z832z4, G932z4, N932z4, U932z4, Ba32z4, Ia32z4, Pa32z4, Wa32z4, Db32z4, Kb32z4;
wire Rb32z4, Yb32z4, Fc32z4, Mc32z4, Tc32z4, Ad32z4, Hd32z4, Od32z4, Vd32z4, Ce32z4;
wire Je32z4, Qe32z4, Xe32z4, Ef32z4, Lf32z4, Sf32z4, Zf32z4, Gg32z4, Ng32z4, Ug32z4;
wire Bh32z4, Ih32z4, Ph32z4, Wh32z4, Di32z4, Ki32z4, Ri32z4, Yi32z4, Fj32z4, Mj32z4;
wire Tj32z4, Ak32z4, Hk32z4, Ok32z4, Vk32z4, Cl32z4, Jl32z4, Ql32z4, Xl32z4, Em32z4;
wire Lm32z4, Sm32z4, Zm32z4, Gn32z4, Nn32z4, Un32z4, Bo32z4, Io32z4, Po32z4, Wo32z4;
wire Dp32z4, Kp32z4, Rp32z4, Yp32z4, Fq32z4, Mq32z4, Tq32z4, Ar32z4, Hr32z4, Or32z4;
wire Vr32z4, Cs32z4, Js32z4, Qs32z4, Xs32z4, Et32z4, Lt32z4, St32z4, Zt32z4, Gu32z4;
wire Nu32z4, Uu32z4, Bv32z4, Iv32z4, Pv32z4, Wv32z4, Dw32z4, Kw32z4, Rw32z4, Yw32z4;
wire Fx32z4, Mx32z4, Tx32z4, Ay32z4, Hy32z4, Oy32z4, Vy32z4, Cz32z4, Jz32z4, Qz32z4;
wire Xz32z4, E042z4, L042z4, S042z4, Z042z4, G142z4, N142z4, U142z4, B242z4, I242z4;
wire P242z4, W242z4, D342z4, K342z4, R342z4, Y342z4, F442z4, M442z4, T442z4, A542z4;
wire H542z4, O542z4, V542z4, C642z4, J642z4, Q642z4, X642z4, E742z4, L742z4, S742z4;
wire Z742z4, G842z4, N842z4, U842z4, B942z4, I942z4, P942z4, W942z4, Da42z4, Ka42z4;
wire Ra42z4, Ya42z4, Fb42z4, Mb42z4, Tb42z4, Ac42z4, Hc42z4, Oc42z4, Vc42z4, Cd42z4;
wire Jd42z4, Qd42z4, Xd42z4, Ee42z4, Le42z4, Se42z4, Ze42z4, Gf42z4, Nf42z4, Uf42z4;
wire Bg42z4, Ig42z4, Pg42z4, Wg42z4, Dh42z4, Kh42z4, Rh42z4, Yh42z4, Fi42z4, Mi42z4;
wire Ti42z4, Aj42z4, Hj42z4, Oj42z4, Vj42z4, Ck42z4, Jk42z4, Qk42z4, Xk42z4, El42z4;
wire Ll42z4, Sl42z4, Zl42z4, Gm42z4, Nm42z4, Um42z4, Bn42z4, In42z4, Pn42z4, Wn42z4;
wire Do42z4, Ko42z4, Ro42z4, Yo42z4, Fp42z4, Mp42z4, Tp42z4, Aq42z4, Hq42z4, Oq42z4;
wire Vq42z4, Cr42z4, Jr42z4, Qr42z4, Xr42z4, Es42z4, Ls42z4, Ss42z4, Zs42z4, Gt42z4;
wire Nt42z4, Ut42z4, Bu42z4, Iu42z4, Pu42z4, Wu42z4, Dv42z4, Kv42z4, Rv42z4, Yv42z4;
wire Fw42z4, Mw42z4, Tw42z4, Ax42z4, Hx42z4, Ox42z4, Vx42z4, Cy42z4, Jy42z4, Qy42z4;
wire Xy42z4, Ez42z4, Lz42z4, Sz42z4, Zz42z4, G052z4, N052z4, U052z4, B152z4, I152z4;
wire P152z4, W152z4, D252z4, K252z4, R252z4, Y252z4, F352z4, M352z4, T352z4, A452z4;
wire H452z4, O452z4, V452z4, C552z4, J552z4, Q552z4, X552z4, E652z4, L652z4, S652z4;
wire Z652z4, G752z4, N752z4, U752z4, B852z4, I852z4, P852z4, W852z4, D952z4, K952z4;
wire R952z4, Y952z4, Fa52z4, Ma52z4, Ta52z4, Ab52z4, Hb52z4, Ob52z4, Vb52z4, Cc52z4;
wire Jc52z4, Qc52z4, Xc52z4, Ed52z4, Ld52z4, Sd52z4, Zd52z4, Ge52z4, Ne52z4, Ue52z4;
wire Bf52z4, If52z4, Pf52z4, Wf52z4, Dg52z4, Kg52z4, Rg52z4, Yg52z4, Fh52z4, Mh52z4;
wire Th52z4, Ai52z4, Hi52z4, Oi52z4, Vi52z4, Cj52z4, Jj52z4, Qj52z4, Xj52z4, Ek52z4;
wire Lk52z4, Sk52z4, Zk52z4, Gl52z4, Nl52z4, Ul52z4, Bm52z4, Im52z4, Pm52z4, Wm52z4;
wire Dn52z4, Kn52z4, Rn52z4, Yn52z4, Fo52z4, Mo52z4, To52z4, Ap52z4, Hp52z4, Op52z4;
wire Vp52z4, Cq52z4, Jq52z4, Qq52z4, Xq52z4, Er52z4, Lr52z4, Sr52z4, Zr52z4, Gs52z4;
wire Ns52z4, Us52z4, Bt52z4, It52z4, Pt52z4, Wt52z4, Du52z4, Ku52z4, Ru52z4, Yu52z4;
wire Fv52z4, Mv52z4, Tv52z4, Aw52z4, Hw52z4, Ow52z4, Vw52z4, Cx52z4, Jx52z4, Qx52z4;
wire Xx52z4, Ey52z4, Ly52z4, Sy52z4, Zy52z4, Gz52z4, Nz52z4, Uz52z4, B062z4, I062z4;
wire P062z4, W062z4, D162z4, K162z4, R162z4, Y162z4, F262z4, M262z4, T262z4, A362z4;
wire H362z4, O362z4, V362z4, C462z4, J462z4, Q462z4, X462z4, E562z4, L562z4, S562z4;
wire Z562z4, G662z4, N662z4, U662z4, B762z4, I762z4, P762z4, W762z4, D862z4, K862z4;
wire R862z4, Y862z4, F962z4, M962z4, T962z4, Aa62z4, Ha62z4, Oa62z4, Va62z4, Cb62z4;
wire Jb62z4, Qb62z4, Xb62z4, Ec62z4, Lc62z4, Sc62z4, Zc62z4, Gd62z4, Nd62z4, Ud62z4;
wire Be62z4, Ie62z4, Pe62z4, We62z4, Df62z4, Kf62z4, Rf62z4, Yf62z4, Fg62z4, Mg62z4;
wire Tg62z4, Ah62z4, Hh62z4, Oh62z4, Vh62z4, Ci62z4, Ji62z4, Qi62z4, Xi62z4, Ej62z4;
wire Lj62z4, Sj62z4, Zj62z4, Gk62z4, Nk62z4, Uk62z4, Bl62z4, Il62z4, Pl62z4, Wl62z4;
wire Dm62z4, Km62z4, Rm62z4, Ym62z4, Fn62z4, Mn62z4, Tn62z4, Ao62z4, Ho62z4, Oo62z4;
wire Vo62z4, Cp62z4, Jp62z4, Qp62z4, Xp62z4, Eq62z4, Lq62z4, Sq62z4, Zq62z4, Gr62z4;
wire Nr62z4, Ur62z4, Bs62z4, Is62z4, Ps62z4, Ws62z4, Dt62z4, Kt62z4, Rt62z4, Yt62z4;
wire Fu62z4, Mu62z4, Tu62z4, Av62z4, Hv62z4, Ov62z4, Vv62z4, Cw62z4, Jw62z4, Qw62z4;
wire Xw62z4, Ex62z4, Lx62z4, Sx62z4, Zx62z4, Gy62z4, Ny62z4, Uy62z4, Bz62z4, Iz62z4;
wire Pz62z4, Wz62z4, D072z4, K072z4, R072z4, Y072z4, F172z4, M172z4, T172z4, A272z4;
wire H272z4, O272z4, V272z4, C372z4, J372z4, Q372z4, X372z4, E472z4, L472z4, S472z4;
wire Z472z4, G572z4, N572z4, U572z4, B672z4, I672z4, P672z4, W672z4, D772z4, K772z4;
wire R772z4, Y772z4, F872z4, M872z4, T872z4, A972z4, H972z4, O972z4, V972z4, Ca72z4;
wire Ja72z4, Qa72z4, Xa72z4, Eb72z4, Lb72z4, Sb72z4, Zb72z4, Gc72z4, Nc72z4, Uc72z4;
wire Bd72z4, Id72z4, Pd72z4, Wd72z4, De72z4, Ke72z4, Re72z4, Ye72z4, Ff72z4, Mf72z4;
wire Tf72z4, Ag72z4, Hg72z4, Og72z4, Vg72z4, Ch72z4, Jh72z4, Qh72z4, Xh72z4, Ei72z4;
wire Li72z4, Si72z4, Zi72z4, Gj72z4, Nj72z4, Uj72z4, Bk72z4, Ik72z4, Pk72z4, Wk72z4;
wire Dl72z4, Kl72z4, Rl72z4, Yl72z4, Fm72z4, Mm72z4, Tm72z4, An72z4, Hn72z4, On72z4;
wire Vn72z4, Co72z4, Jo72z4, Qo72z4, Xo72z4, Ep72z4, Lp72z4, Sp72z4, Zp72z4, Gq72z4;
wire Nq72z4, Uq72z4, Br72z4, Ir72z4, Pr72z4, Wr72z4, Ds72z4, Ks72z4, Rs72z4, Ys72z4;
wire Ft72z4, Mt72z4, Tt72z4, Au72z4, Hu72z4, Ou72z4, Vu72z4, Cv72z4, Jv72z4, Qv72z4;
wire Xv72z4, Ew72z4, Lw72z4, Sw72z4, Zw72z4, Gx72z4, Nx72z4, Ux72z4, By72z4, Iy72z4;
wire Py72z4, Wy72z4, Dz72z4, Kz72z4, Rz72z4, Yz72z4, F082z4, M082z4, T082z4, A182z4;
wire H182z4, O182z4, V182z4, C282z4, J282z4, Q282z4, X282z4, E382z4, L382z4, S382z4;
wire Z382z4, G482z4, N482z4, U482z4, B582z4, I582z4, P582z4, W582z4, D682z4, K682z4;
wire R682z4, Y682z4, F782z4, M782z4, T782z4, A882z4, H882z4, O882z4, V882z4, C982z4;
wire J982z4, Q982z4, X982z4, Ea82z4, La82z4, Sa82z4, Za82z4, Gb82z4, Nb82z4, Ub82z4;
wire Bc82z4, Ic82z4, Pc82z4, Wc82z4, Dd82z4, Kd82z4, Rd82z4, Yd82z4, Fe82z4, Me82z4;
wire Te82z4, Af82z4, Hf82z4, Of82z4, Vf82z4, Cg82z4, Jg82z4, Qg82z4, Xg82z4, Eh82z4;
wire Lh82z4, Sh82z4, Zh82z4, Gi82z4, Ni82z4, Ui82z4, Bj82z4, Ij82z4, Pj82z4, Wj82z4;
wire Dk82z4, Kk82z4, Rk82z4, Yk82z4, Fl82z4, Ml82z4, Tl82z4, Am82z4, Hm82z4, Om82z4;
wire Vm82z4, Cn82z4, Jn82z4, Qn82z4, Xn82z4, Eo82z4, Lo82z4, So82z4, Zo82z4, Gp82z4;
wire Np82z4, Up82z4, Bq82z4, Iq82z4, Pq82z4, Wq82z4, Dr82z4, Kr82z4, Rr82z4, Yr82z4;
wire Fs82z4, Ms82z4, Ts82z4, At82z4, Ht82z4, Ot82z4, Vt82z4, Cu82z4, Ju82z4, Qu82z4;
wire Xu82z4, Ev82z4, Lv82z4, Sv82z4, Zv82z4, Gw82z4, Nw82z4, Uw82z4, Bx82z4, Ix82z4;
wire Px82z4, Wx82z4, Dy82z4, Ky82z4, Ry82z4, Yy82z4, Fz82z4, Mz82z4, Tz82z4, A092z4;
wire H092z4, O092z4, V092z4, C192z4, J192z4, Q192z4, X192z4, E292z4, L292z4, S292z4;
wire Z292z4, G392z4, N392z4, U392z4, B492z4, I492z4, P492z4, W492z4, D592z4, K592z4;
wire R592z4, Y592z4, F692z4, M692z4, T692z4, A792z4, H792z4, O792z4, V792z4, C892z4;
wire J892z4, Q892z4, X892z4, E992z4, L992z4, S992z4, Z992z4, Ga92z4, Na92z4, Ua92z4;
wire Bb92z4, Ib92z4, Pb92z4, Wb92z4, Dc92z4, Kc92z4, Rc92z4, Yc92z4, Fd92z4, Md92z4;
wire Td92z4, Ae92z4, He92z4, Oe92z4, Ve92z4, Cf92z4, Jf92z4, Qf92z4, Xf92z4, Eg92z4;
wire Lg92z4, Sg92z4, Zg92z4, Gh92z4, Nh92z4, Uh92z4, Bi92z4, Ii92z4, Pi92z4, Wi92z4;
wire Dj92z4, Kj92z4, Rj92z4, Yj92z4, Fk92z4, Mk92z4, Tk92z4, Al92z4, Hl92z4, Ol92z4;
wire Vl92z4, Cm92z4, Jm92z4, Qm92z4, Xm92z4, En92z4, Ln92z4, Sn92z4, Zn92z4, Go92z4;
wire No92z4, Uo92z4, Bp92z4, Ip92z4, Pp92z4, Wp92z4, Dq92z4, Kq92z4, Rq92z4, Yq92z4;
wire Fr92z4, Mr92z4, Tr92z4, As92z4, Hs92z4, Os92z4, Vs92z4, Ct92z4, Jt92z4, Qt92z4;
wire Xt92z4, Eu92z4, Lu92z4, Su92z4, Zu92z4, Gv92z4, Nv92z4, Uv92z4, Bw92z4, Iw92z4;
wire Pw92z4, Ww92z4, Dx92z4, Kx92z4, Rx92z4, Yx92z4, Fy92z4, My92z4, Ty92z4, Az92z4;
wire Hz92z4, Oz92z4, Vz92z4, C0a2z4, J0a2z4, Q0a2z4, X0a2z4, E1a2z4, L1a2z4, S1a2z4;
wire Z1a2z4, G2a2z4, N2a2z4, U2a2z4, B3a2z4, I3a2z4, P3a2z4, W3a2z4, D4a2z4, K4a2z4;
wire R4a2z4, Y4a2z4, F5a2z4, M5a2z4, T5a2z4, A6a2z4, H6a2z4, O6a2z4, V6a2z4, C7a2z4;
wire J7a2z4, Q7a2z4, X7a2z4, E8a2z4, L8a2z4, S8a2z4, Z8a2z4, G9a2z4, N9a2z4, U9a2z4;
wire Baa2z4, Iaa2z4, Paa2z4, Waa2z4, Dba2z4, Kba2z4, Rba2z4, Yba2z4, Fca2z4, Mca2z4;
wire Tca2z4, Ada2z4, Hda2z4, Oda2z4, Vda2z4, Cea2z4, Jea2z4, Qea2z4, Xea2z4, Efa2z4;
wire Lfa2z4, Sfa2z4, Zfa2z4, Gga2z4, Nga2z4, Uga2z4, Bha2z4, Iha2z4, Pha2z4, Wha2z4;
wire Dia2z4, Kia2z4, Ria2z4, Yia2z4, Fja2z4, Mja2z4, Tja2z4, Aka2z4, Hka2z4, Oka2z4;
wire Vka2z4, Cla2z4, Jla2z4, Qla2z4, Xla2z4, Ema2z4, Lma2z4, Sma2z4, Zma2z4, Gna2z4;
wire Nna2z4, Una2z4, Boa2z4, Ioa2z4, Poa2z4, Woa2z4, Dpa2z4, Kpa2z4, Rpa2z4, Ypa2z4;
wire Fqa2z4, Mqa2z4, Tqa2z4, Ara2z4, Hra2z4, Ora2z4, Vra2z4, Csa2z4, Jsa2z4, Qsa2z4;
wire Xsa2z4, Eta2z4, Lta2z4, Sta2z4, Zta2z4, Gua2z4, Nua2z4, Uua2z4, Bva2z4, Iva2z4;
wire Pva2z4, Wva2z4, Dwa2z4, Kwa2z4, Rwa2z4, Ywa2z4, Fxa2z4, Mxa2z4, Txa2z4, Aya2z4;
wire Hya2z4, Oya2z4, Vya2z4, Cza2z4, Jza2z4, Qza2z4, Xza2z4, E0b2z4, L0b2z4, S0b2z4;
wire Z0b2z4, G1b2z4, N1b2z4, U1b2z4, B2b2z4, I2b2z4, P2b2z4, W2b2z4, D3b2z4, K3b2z4;
wire R3b2z4, Y3b2z4, F4b2z4, M4b2z4, T4b2z4, A5b2z4, H5b2z4, O5b2z4, V5b2z4, C6b2z4;
wire J6b2z4, Q6b2z4, X6b2z4, E7b2z4, L7b2z4, S7b2z4, Z7b2z4, G8b2z4, N8b2z4, U8b2z4;
wire B9b2z4, I9b2z4, P9b2z4, W9b2z4, Dab2z4, Kab2z4, Rab2z4, Yab2z4, Fbb2z4, Mbb2z4;
wire Tbb2z4, Acb2z4, Hcb2z4, Ocb2z4, Vcb2z4, Cdb2z4, Jdb2z4, Qdb2z4, Xdb2z4, Eeb2z4;
wire Leb2z4, Seb2z4, Zeb2z4, Gfb2z4, Nfb2z4, Ufb2z4, Bgb2z4, Igb2z4, Pgb2z4, Wgb2z4;
wire Dhb2z4, Khb2z4, Rhb2z4, Yhb2z4, Fib2z4, Mib2z4, Tib2z4, Ajb2z4, Hjb2z4, Ojb2z4;
wire Vjb2z4, Ckb2z4, Jkb2z4, Qkb2z4, Xkb2z4, Elb2z4, Llb2z4, Slb2z4, Zlb2z4, Gmb2z4;
wire Nmb2z4, Umb2z4, Bnb2z4, Inb2z4, Pnb2z4, Wnb2z4, Dob2z4, Kob2z4, Rob2z4, Yob2z4;
wire Fpb2z4, Mpb2z4, Tpb2z4, Aqb2z4, Hqb2z4, Oqb2z4, Vqb2z4, Crb2z4, Jrb2z4, Qrb2z4;
wire Xrb2z4, Esb2z4, Lsb2z4, Ssb2z4, Zsb2z4, Gtb2z4, Ntb2z4, Utb2z4, Bub2z4, Iub2z4;
wire Pub2z4, Wub2z4, Dvb2z4, Kvb2z4, Rvb2z4, Yvb2z4, Fwb2z4, Mwb2z4, Twb2z4, Axb2z4;
wire Hxb2z4, Oxb2z4, Vxb2z4, Cyb2z4, Jyb2z4, Qyb2z4, Xyb2z4, Ezb2z4, Lzb2z4, Szb2z4;
wire Zzb2z4, G0c2z4, N0c2z4, U0c2z4, B1c2z4, I1c2z4, P1c2z4, W1c2z4, D2c2z4, K2c2z4;
wire R2c2z4, Y2c2z4, F3c2z4, M3c2z4, T3c2z4, A4c2z4, H4c2z4, O4c2z4, V4c2z4, C5c2z4;
wire J5c2z4, Q5c2z4, X5c2z4, E6c2z4, L6c2z4, S6c2z4, Z6c2z4, G7c2z4, N7c2z4, U7c2z4;
wire B8c2z4, I8c2z4, P8c2z4, W8c2z4, D9c2z4, K9c2z4, R9c2z4, Y9c2z4, Fac2z4, Mac2z4;
wire Tac2z4, Abc2z4, Hbc2z4, Obc2z4, Vbc2z4, Ccc2z4, Jcc2z4, Qcc2z4, Xcc2z4, Edc2z4;
wire Ldc2z4, Sdc2z4, Zdc2z4, Gec2z4, Nec2z4, Uec2z4, Bfc2z4, Ifc2z4, Pfc2z4, Wfc2z4;
wire Dgc2z4, Kgc2z4, Rgc2z4, Ygc2z4, Fhc2z4, Mhc2z4, Thc2z4, Aic2z4, Hic2z4, Oic2z4;
wire Vic2z4, Cjc2z4, Jjc2z4, Qjc2z4, Xjc2z4, Ekc2z4, Lkc2z4, Skc2z4, Zkc2z4, Glc2z4;
wire Nlc2z4, Ulc2z4, Bmc2z4, Imc2z4, Pmc2z4, Wmc2z4, Dnc2z4, Knc2z4, Rnc2z4, Ync2z4;
wire Foc2z4, Moc2z4, Toc2z4, Apc2z4, Hpc2z4, Opc2z4, Vpc2z4, Cqc2z4, Jqc2z4, Qqc2z4;
wire Xqc2z4, Erc2z4, Lrc2z4, Src2z4, Zrc2z4, Gsc2z4, Nsc2z4, Usc2z4, Btc2z4, Itc2z4;
wire Ptc2z4, Wtc2z4, Duc2z4, Kuc2z4, Ruc2z4, Yuc2z4, Fvc2z4, Mvc2z4, Tvc2z4, Awc2z4;
wire Hwc2z4, Owc2z4, Vwc2z4, Cxc2z4, Jxc2z4, Qxc2z4, Xxc2z4, Eyc2z4, Lyc2z4, Syc2z4;
wire Zyc2z4, Gzc2z4, Nzc2z4, Uzc2z4, B0d2z4, I0d2z4, P0d2z4, W0d2z4, D1d2z4, K1d2z4;
wire R1d2z4, Y1d2z4, F2d2z4, M2d2z4, T2d2z4, A3d2z4, H3d2z4, O3d2z4, V3d2z4, C4d2z4;
wire J4d2z4, Q4d2z4, X4d2z4, E5d2z4, L5d2z4, S5d2z4, Z5d2z4, G6d2z4, N6d2z4, U6d2z4;
wire B7d2z4, I7d2z4, P7d2z4, W7d2z4, D8d2z4, K8d2z4, R8d2z4, Y8d2z4, F9d2z4, M9d2z4;
wire T9d2z4, Aad2z4, Had2z4, Oad2z4, Vad2z4, Cbd2z4, Jbd2z4, Qbd2z4, Xbd2z4, Ecd2z4;
wire Lcd2z4, Scd2z4, Zcd2z4, Gdd2z4, Ndd2z4, Udd2z4, Bed2z4, Ied2z4, Ped2z4, Wed2z4;
wire Dfd2z4, Kfd2z4, Rfd2z4, Yfd2z4, Fgd2z4, Mgd2z4, Tgd2z4, Ahd2z4, Hhd2z4, Ohd2z4;
wire Vhd2z4, Cid2z4, Jid2z4, Qid2z4, Xid2z4, Ejd2z4, Ljd2z4, Sjd2z4, Zjd2z4, Gkd2z4;
wire Nkd2z4, Ukd2z4, Bld2z4, Ild2z4, Pld2z4, Wld2z4, Dmd2z4, Kmd2z4, Rmd2z4, Ymd2z4;
wire Fnd2z4, Mnd2z4, Tnd2z4, Aod2z4, Hod2z4, Ood2z4, Vod2z4, Cpd2z4, Jpd2z4, Qpd2z4;
wire Xpd2z4, Eqd2z4, Lqd2z4, Sqd2z4, Zqd2z4, Grd2z4, Nrd2z4, Urd2z4, Bsd2z4, Isd2z4;
wire Psd2z4, Wsd2z4, Dtd2z4, Ktd2z4, Rtd2z4, Ytd2z4, Fud2z4, Mud2z4, Tud2z4, Avd2z4;
wire Hvd2z4, Ovd2z4, Vvd2z4, Cwd2z4, Jwd2z4, Qwd2z4, Xwd2z4, Exd2z4, Lxd2z4, Sxd2z4;
wire Zxd2z4, Gyd2z4, Nyd2z4, Uyd2z4, Bzd2z4, Izd2z4, Pzd2z4, Wzd2z4, D0e2z4, K0e2z4;
wire R0e2z4, Y0e2z4, F1e2z4, M1e2z4, T1e2z4, A2e2z4, H2e2z4, O2e2z4, V2e2z4, C3e2z4;
wire J3e2z4, Q3e2z4, X3e2z4, E4e2z4, L4e2z4, S4e2z4, Z4e2z4, G5e2z4, N5e2z4, U5e2z4;
wire B6e2z4, I6e2z4, P6e2z4, W6e2z4, D7e2z4, K7e2z4, R7e2z4, Y7e2z4, F8e2z4, M8e2z4;
wire T8e2z4, A9e2z4, H9e2z4, O9e2z4, V9e2z4, Cae2z4, Jae2z4, Qae2z4, Xae2z4, Ebe2z4;
wire Lbe2z4, Sbe2z4, Zbe2z4, Gce2z4, Nce2z4, Uce2z4, Bde2z4, Ide2z4, Pde2z4, Wde2z4;
wire Dee2z4, Kee2z4, Ree2z4, Yee2z4, Ffe2z4, Mfe2z4, Tfe2z4, Age2z4, Hge2z4, Oge2z4;
wire Vge2z4, Che2z4, Jhe2z4, Qhe2z4, Xhe2z4, Eie2z4, Lie2z4, Sie2z4, Zie2z4, Gje2z4;
wire Nje2z4, Uje2z4, Bke2z4, Ike2z4, Pke2z4, Wke2z4, Dle2z4, Kle2z4, Rle2z4, Yle2z4;
wire Fme2z4, Mme2z4, Tme2z4, Ane2z4, Hne2z4, One2z4, Vne2z4, Coe2z4, Joe2z4, Qoe2z4;
wire Xoe2z4, Epe2z4, Lpe2z4, Spe2z4, Zpe2z4, Gqe2z4, Nqe2z4, Uqe2z4, Bre2z4, Ire2z4;
wire Pre2z4, Wre2z4, Dse2z4, Kse2z4, Rse2z4, Yse2z4, Fte2z4, Mte2z4, Tte2z4, Aue2z4;
wire Hue2z4, Oue2z4, Vue2z4, Cve2z4, Jve2z4, Qve2z4, Xve2z4, Ewe2z4, Lwe2z4, Swe2z4;
wire Zwe2z4, Gxe2z4, Nxe2z4, Uxe2z4, Bye2z4, Iye2z4, Pye2z4, Wye2z4, Dze2z4, Kze2z4;
wire Rze2z4, Yze2z4, F0f2z4, M0f2z4, T0f2z4, A1f2z4, H1f2z4, O1f2z4, V1f2z4, C2f2z4;
wire J2f2z4, Q2f2z4, X2f2z4, E3f2z4, L3f2z4, S3f2z4, Z3f2z4, G4f2z4, N4f2z4, U4f2z4;
wire B5f2z4, I5f2z4, P5f2z4, W5f2z4, D6f2z4, K6f2z4, R6f2z4, Y6f2z4, F7f2z4, M7f2z4;
wire T7f2z4, A8f2z4, H8f2z4, O8f2z4, V8f2z4, C9f2z4, J9f2z4, Q9f2z4, X9f2z4, Eaf2z4;
wire Laf2z4, Saf2z4, Zaf2z4, Gbf2z4, Nbf2z4, Ubf2z4, Bcf2z4, Icf2z4, Pcf2z4, Wcf2z4;
wire Ddf2z4, Kdf2z4, Rdf2z4, Ydf2z4, Fef2z4, Mef2z4, Tef2z4, Aff2z4, Hff2z4, Off2z4;
wire Vff2z4, Cgf2z4, Jgf2z4, Qgf2z4, Xgf2z4, Ehf2z4, Lhf2z4, Shf2z4, Zhf2z4, Gif2z4;
wire Nif2z4, Uif2z4, Bjf2z4, Ijf2z4, Pjf2z4, Wjf2z4, Dkf2z4, Kkf2z4, Rkf2z4, Ykf2z4;
wire Flf2z4, Mlf2z4, Tlf2z4, Amf2z4, Hmf2z4, Omf2z4, Vmf2z4, Cnf2z4, Jnf2z4, Qnf2z4;
wire Xnf2z4, Eof2z4, Lof2z4, Sof2z4, Zof2z4, Gpf2z4, Npf2z4, Upf2z4, Bqf2z4, Iqf2z4;
wire Pqf2z4, Wqf2z4, Drf2z4, Krf2z4, Rrf2z4, Yrf2z4, Fsf2z4, Msf2z4, Tsf2z4, Atf2z4;
wire Htf2z4, Otf2z4, Vtf2z4, Cuf2z4, Juf2z4, Quf2z4, Xuf2z4, Evf2z4, Lvf2z4, Svf2z4;
wire Zvf2z4, Gwf2z4, Nwf2z4, Uwf2z4, Bxf2z4, Ixf2z4, Pxf2z4, Wxf2z4, Dyf2z4, Kyf2z4;
wire Ryf2z4, Yyf2z4, Fzf2z4, Mzf2z4, Tzf2z4, A0g2z4, H0g2z4, O0g2z4, V0g2z4, C1g2z4;
wire J1g2z4, Q1g2z4, X1g2z4, E2g2z4, L2g2z4, S2g2z4, Z2g2z4, G3g2z4, N3g2z4, U3g2z4;
wire B4g2z4, I4g2z4, P4g2z4, W4g2z4, D5g2z4, K5g2z4, R5g2z4, Y5g2z4, F6g2z4, M6g2z4;
wire T6g2z4, A7g2z4, H7g2z4, O7g2z4, V7g2z4, C8g2z4, J8g2z4, Q8g2z4, X8g2z4, E9g2z4;
wire L9g2z4, S9g2z4, Z9g2z4, Gag2z4, Nag2z4, Uag2z4, Bbg2z4, Ibg2z4, Pbg2z4, Wbg2z4;
wire Dcg2z4, Kcg2z4, Rcg2z4, Ycg2z4, Fdg2z4, Mdg2z4, Tdg2z4, Aeg2z4, Heg2z4, Oeg2z4;
wire Veg2z4, Cfg2z4, Jfg2z4, Qfg2z4, Xfg2z4, Egg2z4, Lgg2z4, Sgg2z4, Zgg2z4, Ghg2z4;
wire Nhg2z4, Uhg2z4, Big2z4, Iig2z4, Pig2z4, Wig2z4, Djg2z4, Kjg2z4, Rjg2z4, Yjg2z4;
wire Fkg2z4, Mkg2z4, Tkg2z4, Alg2z4, Hlg2z4, Olg2z4, Vlg2z4, Cmg2z4, Jmg2z4, Qmg2z4;
wire Xmg2z4, Eng2z4, Lng2z4, Sng2z4, Zng2z4, Gog2z4, Nog2z4, Uog2z4, Bpg2z4, Ipg2z4;
wire Ppg2z4, Wpg2z4, Dqg2z4, Kqg2z4, Rqg2z4, Yqg2z4, Frg2z4, Mrg2z4, Trg2z4, Asg2z4;
wire Hsg2z4, Osg2z4, Vsg2z4, Ctg2z4, Jtg2z4, Qtg2z4, Xtg2z4, Eug2z4, Lug2z4, Sug2z4;
wire Zug2z4, Gvg2z4, Nvg2z4, Uvg2z4, Bwg2z4, Iwg2z4, Pwg2z4, Wwg2z4, Dxg2z4, Kxg2z4;
wire Rxg2z4, Yxg2z4, Fyg2z4, Myg2z4, Tyg2z4, Azg2z4, Hzg2z4, Ozg2z4, Vzg2z4, C0h2z4;
wire J0h2z4, Q0h2z4, X0h2z4, E1h2z4, L1h2z4, S1h2z4, Z1h2z4, G2h2z4, N2h2z4, U2h2z4;
wire B3h2z4, I3h2z4, P3h2z4, W3h2z4, D4h2z4, K4h2z4, R4h2z4, Y4h2z4, F5h2z4, M5h2z4;
wire T5h2z4, A6h2z4, H6h2z4, O6h2z4, V6h2z4, C7h2z4, J7h2z4, Q7h2z4, X7h2z4, E8h2z4;
wire L8h2z4, S8h2z4, Z8h2z4, G9h2z4, N9h2z4, U9h2z4, Bah2z4, Iah2z4, Pah2z4, Wah2z4;
wire Dbh2z4, Kbh2z4, Rbh2z4, Ybh2z4, Fch2z4, Mch2z4, Tch2z4, Adh2z4, Hdh2z4, Odh2z4;
wire Vdh2z4, Ceh2z4, Jeh2z4, Qeh2z4, Xeh2z4, Efh2z4, Lfh2z4, Sfh2z4, Zfh2z4, Ggh2z4;
wire Ngh2z4, Ugh2z4, Bhh2z4, Ihh2z4, Phh2z4, Whh2z4, Dih2z4, Kih2z4, Rih2z4, Yih2z4;
wire Fjh2z4, Mjh2z4;
wire [3:0] Tjh2z4;
wire [30:2] Ykh2z4;
wire [31:0] Dmh2z4;
wire [8:1] Enh2z4;
wire [30:0] Roh2z4;
wire [1:0] Zph2z4;
wire [23:0] Irh2z4;
wire [1:0] Psh2z4;
wire [1:0] Uth2z4;
wire [31:0] Zuh2z4;
wire [23:0] Iwh2z4;
wire [1:0] Txh2z4;
wire [23:0] Czh2z4;
wire [15:0] L0i2z4;
wire [15:0] T1i2z4;
wire [15:0] D3i2z4;
wire N4i2z4, L5i2z4;
reg J6i2z4, Z7i2z4, H9i2z4, Wai2z4, Gci2z4, Pdi2z4, Zei2z4, Igi2z4, Rhi2z4, Gji2z4;
reg Tki2z4, Emi2z4, Rni2z4, Fpi2z4, Uqi2z4, Isi2z4, Xti2z4, Mvi2z4, Ywi2z4, Kyi2z4;
reg Yzi2z4, M1j2z4, X2j2z4, M4j2z4, B6j2z4, Q7j2z4, F9j2z4, Uaj2z4, Fcj2z4, Qdj2z4;
reg Ffj2z4, Sgj2z4, Fij2z4, Sjj2z4, Glj2z4, Vmj2z4, Koj2z4, Zpj2z4, Orj2z4, Dtj2z4;
reg Ruj2z4, Fwj2z4, Txj2z4, Hzj2z4, V0k2z4, K2k2z4, Z3k2z4, O5k2z4, D7k2z4, S8k2z4;
reg Hak2z4, Wbk2z4, Idk2z4, Rek2z4, Ggk2z4, Vhk2z4, Kjk2z4, Zkk2z4, Omk2z4, Aok2z4;
reg Npk2z4, Ark2z4, Nsk2z4, Auk2z4, Svk2z4, Gxk2z4, Xyk2z4, J0l2z4, V1l2z4, K3l2z4;
reg Z4l2z4, Q6l2z4, H8l2z4, Y9l2z4, Pbl2z4, Edl2z4, Tel2z4, Igl2z4, Xhl2z4, Mjl2z4;
reg Cll2z4, Qml2z4, Eol2z4, Spl2z4, Grl2z4, Usl2z4, Lul2z4, Dwl2z4, Rxl2z4, Fzl2z4;
reg T0m2z4, H2m2z4, V3m2z4, J5m2z4, X6m2z4, L8m2z4, Cam2z4, Nbm2z4, Bdm2z4, Qem2z4;
reg Fgm2z4, Thm2z4, Ejm2z4, Skm2z4, Gmm2z4, Unm2z4, Ipm2z4, Wqm2z4, Ksm2z4, Ytm2z4;
reg Mvm2z4, Axm2z4, Rym2z4, J0n2z4, Y1n2z4, N3n2z4, C5n2z4, R6n2z4, G8n2z4, X9n2z4;
reg Lbn2z4, Zcn2z4, Nen2z4, Yfn2z4, Mhn2z4, Ajn2z4, Okn2z4, Cmn2z4, Qnn2z4, Ipn2z4;
reg Arn2z4, Psn2z4, Eun2z4, Tvn2z4, Ixn2z4, Xyn2z4, O0o2z4, F2o2z4, V3o2z4, J5o2z4;
reg Y6o2z4, N8o2z4, Cao2z4, Rbo2z4, Gdo2z4, Xeo2z4, Ogo2z4, Fio2z4, Ujo2z4, Jlo2z4;
reg Ymo2z4, Noo2z4, Cqo2z4, Rro2z4, Gto2z4, Vuo2z4, Kwo2z4, Zxo2z4, Ozo2z4, D1p2z4;
reg S2p2z4, H4p2z4, W5p2z4, L7p2z4, A9p2z4, Pap2z4, Ecp2z4, Tdp2z4, Efp2z4, Sgp2z4;
reg Gip2z4, Ujp2z4, Ilp2z4, Wmp2z4, Kop2z4, Aqp2z4, Qrp2z4, Gtp2z4, Uup2z4, Iwp2z4;
reg Wxp2z4, Mzp2z4, B1q2z4, Q2q2z4, F4q2z4, U5q2z4, J7q2z4, Y8q2z4, Naq2z4, Ccq2z4;
reg Rdq2z4, Gfq2z4, Vgq2z4, Kiq2z4, Zjq2z4, Llq2z4, Anq2z4, Poq2z4, Eqq2z4, Trq2z4;
reg Etq2z4, Wuq2z4, Owq2z4, Cyq2z4, Qzq2z4, E1r2z4, S2r2z4, G4r2z4, U5r2z4, I7r2z4;
reg W8r2z4, Oar2z4, Gcr2z4, Vdr2z4, Kfr2z4, Zgr2z4, Oir2z4, Dkr2z4, Slr2z4, Hnr2z4;
reg Wor2z4, Lqr2z4, Asr2z4, Otr2z4, Cvr2z4, Qwr2z4, Eyr2z4, Szr2z4, G1s2z4, U2s2z4;
reg I4s2z4, W5s2z4, K7s2z4, Z8s2z4, Oas2z4, Dcs2z4, Rds2z4, Ffs2z4, Vgs2z4, Mis2z4;
reg Dks2z4, Uls2z4, Lns2z4, Cps2z4, Tqs2z4, Kss2z4, Bus2z4, Svs2z4, Jxs2z4, Azs2z4;
reg R0t2z4, I2t2z4, A4t2z4, O5t2z4, Y6t2z4, L8t2z4, Y9t2z4, Mbt2z4, Adt2z4, Pet2z4;
reg Cgt2z4, Rht2z4, Gjt2z4, Ukt2z4, Imt2z4, Wnt2z4, Lpt2z4, Art2z4, Pst2z4, Eut2z4;
reg Tvt2z4, Ixt2z4, Wyt2z4, K0u2z4, Y1u2z4, M3u2z4, B5u2z4, Q6u2z4, F8u2z4, U9u2z4;
reg Jbu2z4, Ycu2z4, Neu2z4, Cgu2z4, Rhu2z4, Gju2z4, Uku2z4, Imu2z4, Wnu2z4, Lpu2z4;
reg Aru2z4, Psu2z4, Duu2z4, Rvu2z4, Fxu2z4, Uyu2z4, J0v2z4, Y1v2z4, N3v2z4, C5v2z4;
reg R6v2z4, F8v2z4, T9v2z4, Hbv2z4, Vcv2z4, Kev2z4, Zfv2z4, Ohv2z4, Djv2z4, Skv2z4;
reg Hmv2z4, Wnv2z4, Lpv2z4, Arv2z4, Psv2z4, Duv2z4, Rvv2z4, Fxv2z4, Uyv2z4, G0w2z4;
reg R1w2z4, C3w2z4, S4w2z4, I6w2z4, U7w2z4, G9w2z4, Vaw2z4, Jcw2z4, Ydw2z4, Mfw2z4;
reg Ahw2z4, Oiw2z4, Ckw2z4, Qlw2z4, Enw2z4, Sow2z4, Gqw2z4, Urw2z4, Itw2z4, Xuw2z4;
reg Mww2z4, Byw2z4, Qzw2z4, F1x2z4, U2x2z4, J4x2z4, U5x2z4, G7x2z4, R8x2z4, Cax2z4;
reg Nbx2z4, Ycx2z4, Jex2z4, Ufx2z4, Fhx2z4, Rix2z4, Dkx2z4, Plx2z4, Bnx2z4, Nox2z4;
reg Zpx2z4, Lrx2z4, Xsx2z4, Jux2z4, Vvx2z4, Hxx2z4, Tyx2z4, F0y2z4, T1y2z4, I3y2z4;
reg W4y2z4, K6y2z4, Y7y2z4, M9y2z4, Bby2z4, Qcy2z4, Fey2z4, Ufy2z4, Jhy2z4, Viy2z4;
reg Jky2z4, Xly2z4, Lny2z4, Zoy2z4, Nqy2z4, Bsy2z4, Pty2z4, Dvy2z4, Swy2z4, Hyy2z4;
reg Wzy2z4, K1z2z4, C3z2z4, U4z2z4, I6z2z4, W7z2z4, K9z2z4, Yaz2z4, Mcz2z4, Aez2z4;
reg Pfz2z4, Ehz2z4, Tiz2z4, Ikz2z4, Wlz2z4, Knz2z4, Yoz2z4, Nqz2z4, Csz2z4, Rtz2z4;
reg Fvz2z4, Twz2z4, Hyz2z4, Vzz2z4, K103z4, Z203z4, O403z4, D603z4, S703z4, H903z4;
reg Wa03z4, Kc03z4, Yd03z4, Nf03z4, Ch03z4, Qi03z4, Ek03z4, Sl03z4, Hn03z4, Wo03z4;
reg Lq03z4, Zr03z4, Nt03z4, Bv03z4, Pw03z4, Ey03z4, Tz03z4, I113z4, X213z4, M413z4;
reg B613z4, Q713z4, E913z4, Sa13z4, Hc13z4, Wd13z4, Kf13z4, Yg13z4, Mi13z4, Bk13z4;
reg Ql13z4, Fn13z4, Uo13z4, Jq13z4, Yr13z4, Mt13z4, Av13z4, Ow13z4, Cy13z4, Rz13z4;
reg G123z4, V223z4, K423z4, Z523z4, O723z4, D923z4, Sa23z4, Hc23z4, Wd23z4, Kf23z4;
reg Yg23z4, Mi23z4, Bk23z4, Ql23z4, Fn23z4, To23z4, Hq23z4, Vr23z4, Kt23z4, Zu23z4;
reg Ow23z4, Dy23z4, Sz23z4, H133z4, V233z4, J433z4, X533z4, L733z4, A933z4, Pa33z4;
reg Ec33z4, Td33z4, If33z4, Xg33z4, Mi33z4, Bk33z4, Ql33z4, Fn33z4, To33z4, Hq33z4;
reg Vr33z4, Kt33z4, Zu33z4, Ow33z4, Cy33z4, Qz33z4, E143z4, T243z4, I443z4, X543z4;
reg M743z4, B943z4, Qa43z4, Ec43z4, Sd43z4, Gf43z4, Ug43z4, Ji43z4, Yj43z4, Nl43z4;
reg Cn43z4, Ro43z4, Gq43z4, Vr43z4, Kt43z4, Zu43z4, Ow43z4, Cy43z4, Qz43z4, E153z4;
reg T253z4, I453z4, X553z4, L753z4, Z853z4, Na53z4, Cc53z4, Rd53z4, Gf53z4, Vg53z4;
reg Ki53z4, Zj53z4, Nl53z4, Bn53z4, Po53z4, Dq53z4, Sr53z4, Ht53z4, Wu53z4, Lw53z4;
reg Ay53z4, Pz53z4, E163z4, T263z4, I463z4, X563z4, L763z4, Z863z4, Na63z4, Cc63z4;
reg Rd63z4, Gf63z4, Ug63z4, Ii63z4, Wj63z4, Ll63z4, An63z4, Po63z4, Eq63z4, Tr63z4;
reg It63z4, Wu63z4, Kw63z4, Yx63z4, Mz63z4, B173z4, Q273z4, F473z4, U573z4, J773z4;
reg Y873z4, Na73z4, Cc73z4, Rd73z4, Gf73z4, Ug73z4, Ii73z4, Wj73z4, Ll73z4, An73z4;
reg Po73z4, Dq73z4, Rr73z4, Ft73z4, Uu73z4, Jw73z4, Yx73z4, Nz73z4, C183z4, R283z4;
reg F483z4, T583z4, H783z4, V883z4, Ka83z4, Zb83z4, Od83z4, Df83z4, Sg83z4, Hi83z4;
reg Wj83z4, Ll83z4, An83z4, Po83z4, Dq83z4, Rr83z4, Ft83z4, Uu83z4, Jw83z4, Yx83z4;
reg Nz83z4, C193z4, R293z4, G493z4, U593z4, I793z4, W893z4, Ka93z4, Yb93z4, Md93z4;
reg Bf93z4, Qg93z4, Fi93z4, Uj93z4, Jl93z4, Ym93z4, No93z4, Cq93z4, Rr93z4, Gt93z4;
reg Vu93z4, Jw93z4, Xx93z4, Lz93z4, B1a3z4, P2a3z4, D4a3z4, U5a3z4, L7a3z4, C9a3z4;
reg Taa3z4, Jca3z4, Aea3z4, Qfa3z4, Gha3z4, Wia3z4, Mka3z4, Cma3z4, Tna3z4, Jpa3z4;
reg Ara3z4, Rsa3z4, Iua3z4, Zva3z4, Qxa3z4, Gza3z4, W0b3z4, M2b3z4, C4b3z4, S5b3z4;
reg J7b3z4, Z8b3z4, Pab3z4, Gcb3z4, Xdb3z4, Nfb3z4, Dhb3z4, Tib3z4, Kkb3z4, Bmb3z4;
reg Rnb3z4, Ipb3z4, Zqb3z4, Qsb3z4, Hub3z4, Yvb3z4, Pxb3z4, Gzb3z4, X0c3z4, O2c3z4;
reg F4c3z4, W5c3z4, N7c3z4, E9c3z4, Vac3z4, Mcc3z4, Bec3z4, Qfc3z4, Fhc3z4, Uic3z4;
reg Jkc3z4, Ylc3z4, Nnc3z4, Dpc3z4, Tqc3z4, Jsc3z4, Ztc3z4, Ovc3z4, Cxc3z4, Qyc3z4;
reg E0d3z4, T1d3z4, H3d3z4, V4d3z4, G6d3z4, T7d3z4, J9d3z4, Zad3z4, Pcd3z4, Fed3z4;
reg Vfd3z4, Lhd3z4, Bjd3z4, Rkd3z4, Gmd3z4, Snd3z4, Hpd3z4, Wqd3z4, Lsd3z4, Aud3z4;
reg Pvd3z4, Exd3z4, Tyd3z4, I0e3z4, X1e3z4, M3e3z4, B5e3z4, Q6e3z4, F8e3z4, U9e3z4;
reg Ibe3z4, Wce3z4, Lee3z4, Bge3z4, She3z4, Jje3z4, Ble3z4, Tme3z4, Foe3z4, Rpe3z4;
reg Fre3z4, Tse3z4, Hue3z4, Vve3z4, Kxe3z4, Aze3z4, Q0f3z4, H2f3z4, W3f3z4, M5f3z4;
reg C7f3z4, T8f3z4, Kaf3z4, Wbf3z4, Ldf3z4, Aff3z4, Pgf3z4, Eif3z4, Tjf3z4, Ilf3z4;
reg Xmf3z4, Mof3z4, Bqf3z4, Qrf3z4, Ftf3z4, Uuf3z4, Jwf3z4, Vxf3z4, Kzf3z4, Z0g3z4;
reg O2g3z4, D4g3z4, T5g3z4, K7g3z4, B9g3z4, Nag3z4, Ccg3z4, Rdg3z4, Gfg3z4, Vgg3z4;
reg Kig3z4, Zjg3z4, Olg3z4, Dng3z4, Sog3z4, Hqg3z4, Wrg3z4, Ltg3z4, Avg3z4, Pwg3z4;
reg Eyg3z4, Tzg3z4, I1h3z4, Z2h3z4, Q4h3z4, I6h3z4, A8h3z4, P9h3z4, Ebh3z4, Tch3z4;
reg Ieh3z4, Zfh3z4, Ohh3z4, Djh3z4, Skh3z4, Hmh3z4, Wnh3z4, Lph3z4, Arh3z4, Psh3z4;
reg Euh3z4, Tvh3z4, Ixh3z4, Xyh3z4, M0i3z4, B2i3z4, S3i3z4, J5i3z4, Y6i3z4, N8i3z4;
reg Cai3z4, Rbi3z4, Ddi3z4, Uei3z4, Lgi3z4, Aii3z4, Qji3z4, Fli3z4, Umi3z4, Joi3z4;
reg Ypi3z4;
wire [33:0] Pri3z4;
wire [33:0] Fti3z4;

assign hprot_o[1] = 1'b1;
assign hburst_o[2] = 1'b0;
assign hburst_o[1] = 1'b0;
assign hburst_o[0] = 1'b0;
assign hmastlock_o = 1'b0;
assign hsize_o[2] = 1'b0;
assign htrans_o[0] = 1'b0;
assign Xahvx4 = J6i2z4;
assign vis_tbit_o = Z7i2z4;
assign Sh9vx4 = H9i2z4;
assign Dw8vx4 = Wai2z4;
assign vis_apsr_o[3] = Gci2z4;
assign O8gvx4 = Pdi2z4;
assign vis_apsr_o[1] = Zei2z4;
assign vis_apsr_o[2] = Igi2z4;
assign S4evx4 = Rhi2z4;
assign Ih8vx4 = Gji2z4;
assign Cn8vx4 = Tki2z4;
assign Whgvx4 = Emi2z4;
assign Tjh2z4[3] = Rni2z4;
assign vis_r7_o[23] = Fpi2z4;
assign Psh2z4[1] = Uqi2z4;
assign vis_r7_o[31] = Isi2z4;
assign vis_r0_o[31] = Xti2z4;
assign Aygvx4 = Mvi2z4;
assign Eqgvx4 = Ywi2z4;
assign Hnevx4 = Kyi2z4;
assign Uz8vx4 = Yzi2z4;
assign O7evx4 = M1j2z4;
assign vis_msp_o[29] = X2j2z4;
assign vis_msp_o[21] = M4j2z4;
assign Tudvx4 = B6j2z4;
assign Ewdvx4 = Q7j2z4;
assign vis_r7_o[24] = F9j2z4;
assign vis_ipsr_o[2] = Uaj2z4;
assign vis_pc_o[0] = Fcj2z4;
assign Ho8vx4 = Qdj2z4;
assign Nggvx4 = Ffj2z4;
assign Efgvx4 = Sgj2z4;
assign Mcgvx4 = Fij2z4;
assign Tjh2z4[0] = Sjj2z4;
assign vis_r5_o[31] = Glj2z4;
assign vis_r5_o[24] = Vmj2z4;
assign vis_r1_o[31] = Koj2z4;
assign vis_r1_o[24] = Zpj2z4;
assign vis_r1_o[23] = Orj2z4;
assign vis_r5_o[1] = Dtj2z4;
assign vis_r7_o[1] = Ruj2z4;
assign vis_r1_o[1] = Fwj2z4;
assign vis_r0_o[1] = Txj2z4;
assign R3hvx4 = Hzj2z4;
assign vis_r1_o[26] = V0k2z4;
assign vis_r5_o[26] = K2k2z4;
assign vis_r7_o[26] = Z3k2z4;
assign vis_msp_o[24] = O5k2z4;
assign vis_psp_o[24] = D7k2z4;
assign Azdvx4 = S8k2z4;
assign L0evx4 = Hak2z4;
assign Qsgvx4 = Wbk2z4;
assign vis_apsr_o[0] = Idk2z4;
assign vis_msp_o[26] = Rek2z4;
assign vis_r5_o[28] = Ggk2z4;
assign vis_r7_o[28] = Vhk2z4;
assign vis_r1_o[28] = Kjk2z4;
assign vis_r0_o[28] = Zkk2z4;
assign vis_pc_o[29] = Omk2z4;
assign Dbgvx4 = Aok2z4;
assign U9gvx4 = Npk2z4;
assign Z6gvx4 = Ark2z4;
assign Vdgvx4 = Nsk2z4;
assign Su9vx4 = Auk2z4;
assign Xq8vx4 = Svk2z4;
assign T1i2z4[0] = Gxk2z4;
assign vis_pc_o[23] = Xyk2z4;
assign vis_pc_o[30] = J0l2z4;
assign D6evx4 = V1l2z4;
assign Mf8vx4 = K3l2z4;
assign Zuh2z4[13] = Z4l2z4;
assign Zuh2z4[14] = Q6l2z4;
assign Zuh2z4[15] = H8l2z4;
assign T1i2z4[9] = Y9l2z4;
assign vis_r1_o[25] = Pbl2z4;
assign vis_r5_o[25] = Edl2z4;
assign vis_r7_o[25] = Tel2z4;
assign vis_msp_o[23] = Igl2z4;
assign vis_psp_o[23] = Xhl2z4;
assign B5hvx4 = Mjl2z4;
assign vis_msp_o[5] = Cll2z4;
assign vis_r5_o[7] = Qml2z4;
assign vis_r7_o[7] = Eol2z4;
assign vis_r1_o[7] = Spl2z4;
assign vis_r0_o[7] = Grl2z4;
assign Zuh2z4[11] = Usl2z4;
assign T1i2z4[15] = Lul2z4;
assign Roevx4 = Dwl2z4;
assign B19vx4 = Rxl2z4;
assign Ml9vx4 = Fzl2z4;
assign vis_r1_o[3] = T0m2z4;
assign vis_r5_o[3] = H2m2z4;
assign vis_r7_o[3] = V3m2z4;
assign vis_msp_o[1] = J5m2z4;
assign vis_psp_o[1] = X6m2z4;
assign Czh2z4[19] = L8m2z4;
assign vis_ipsr_o[3] = Cam2z4;
assign Xlevx4 = Nbm2z4;
assign K5fvx4 = Bdm2z4;
assign Kg9vx4 = Qem2z4;
assign Tjh2z4[1] = Fgm2z4;
assign vis_primask_o = Thm2z4;
assign vis_r5_o[0] = Ejm2z4;
assign vis_r7_o[0] = Skm2z4;
assign vis_r1_o[0] = Gmm2z4;
assign vis_r0_o[0] = Unm2z4;
assign vis_r1_o[6] = Ipm2z4;
assign vis_r5_o[6] = Wqm2z4;
assign vis_r7_o[6] = Ksm2z4;
assign vis_msp_o[4] = Ytm2z4;
assign vis_psp_o[4] = Mvm2z4;
assign Zuh2z4[10] = Axm2z4;
assign T1i2z4[14] = Rym2z4;
assign vis_r1_o[22] = J0n2z4;
assign vis_r5_o[22] = Y1n2z4;
assign vis_r7_o[22] = N3n2z4;
assign vis_msp_o[20] = C5n2z4;
assign vis_psp_o[20] = R6n2z4;
assign Zuh2z4[12] = G8n2z4;
assign Psh2z4[0] = X9n2z4;
assign Bqevx4 = Lbn2z4;
assign Qm9vx4 = Zcn2z4;
assign vis_control_o = Nen2z4;
assign vis_r1_o[2] = Yfn2z4;
assign vis_r5_o[2] = Mhn2z4;
assign vis_r7_o[2] = Ajn2z4;
assign vis_msp_o[0] = Okn2z4;
assign vis_psp_o[0] = Cmn2z4;
assign D3i2z4[10] = Qnn2z4;
assign T1i2z4[10] = Ipn2z4;
assign vis_r1_o[18] = Arn2z4;
assign vis_r5_o[18] = Psn2z4;
assign vis_r7_o[18] = Eun2z4;
assign vis_msp_o[16] = Tvn2z4;
assign vis_psp_o[16] = Ixn2z4;
assign Czh2z4[18] = Xyn2z4;
assign Irh2z4[18] = O0o2z4;
assign Irh2z4[0] = F2o2z4;
assign Izgvx4 = V3o2z4;
assign vis_r1_o[16] = J5o2z4;
assign vis_r5_o[16] = Y6o2z4;
assign vis_r7_o[16] = N8o2z4;
assign vis_msp_o[14] = Cao2z4;
assign vis_psp_o[14] = Rbo2z4;
assign Czh2z4[16] = Gdo2z4;
assign Irh2z4[16] = Xeo2z4;
assign Irh2z4[21] = Ogo2z4;
assign vis_r1_o[29] = Fio2z4;
assign vis_r5_o[29] = Ujo2z4;
assign vis_r7_o[29] = Jlo2z4;
assign vis_msp_o[27] = Ymo2z4;
assign vis_psp_o[27] = Noo2z4;
assign H3evx4 = Cqo2z4;
assign vis_r1_o[30] = Rro2z4;
assign vis_r5_o[30] = Gto2z4;
assign vis_r7_o[30] = Vuo2z4;
assign vis_r1_o[17] = Kwo2z4;
assign vis_r5_o[17] = Zxo2z4;
assign vis_r7_o[17] = Ozo2z4;
assign vis_msp_o[15] = D1p2z4;
assign vis_psp_o[15] = S2p2z4;
assign Fmdvx4 = H4p2z4;
assign Qndvx4 = W5p2z4;
assign Bpdvx4 = L7p2z4;
assign vis_r1_o[19] = A9p2z4;
assign vis_r5_o[19] = Pap2z4;
assign vis_r7_o[19] = Ecp2z4;
assign vis_ipsr_o[5] = Tdp2z4;
assign I5dvx4 = Efp2z4;
assign vis_r1_o[5] = Sgp2z4;
assign vis_r5_o[5] = Gip2z4;
assign vis_r7_o[5] = Ujp2z4;
assign vis_msp_o[3] = Ilp2z4;
assign vis_psp_o[3] = Wmp2z4;
assign L9hvx4 = Kop2z4;
assign Txh2z4[0] = Aqp2z4;
assign Txh2z4[1] = Qrp2z4;
assign Lrevx4 = Gtp2z4;
assign Un9vx4 = Uup2z4;
assign Kycvx4 = Iwp2z4;
assign Zph2z4[1] = Wxp2z4;
assign vis_r1_o[14] = Mzp2z4;
assign vis_r5_o[14] = B1q2z4;
assign vis_r7_o[14] = Q2q2z4;
assign vis_msp_o[12] = F4q2z4;
assign vis_psp_o[12] = U5q2z4;
assign Yhdvx4 = J7q2z4;
assign Jjdvx4 = Y8q2z4;
assign vis_r1_o[15] = Naq2z4;
assign vis_r5_o[15] = Ccq2z4;
assign vis_r7_o[15] = Rdq2z4;
assign vis_r1_o[27] = Gfq2z4;
assign vis_r5_o[27] = Vgq2z4;
assign vis_r7_o[27] = Kiq2z4;
assign vis_pc_o[18] = Zjq2z4;
assign Xrdvx4 = Llq2z4;
assign vis_r1_o[21] = Anq2z4;
assign vis_r5_o[21] = Poq2z4;
assign vis_r7_o[21] = Eqq2z4;
assign vis_ipsr_o[4] = Trq2z4;
assign D3i2z4[13] = Etq2z4;
assign T1i2z4[13] = Wuq2z4;
assign Vsevx4 = Owq2z4;
assign Yo9vx4 = Cyq2z4;
assign Ik9vx4 = Qzq2z4;
assign vis_r1_o[4] = E1r2z4;
assign vis_r5_o[4] = S2r2z4;
assign vis_r7_o[4] = G4r2z4;
assign vis_msp_o[2] = U5r2z4;
assign vis_psp_o[2] = I7r2z4;
assign D3i2z4[12] = W8r2z4;
assign T1i2z4[12] = Oar2z4;
assign vis_r1_o[12] = Gcr2z4;
assign vis_r5_o[12] = Vdr2z4;
assign vis_r7_o[12] = Kfr2z4;
assign vis_msp_o[10] = Zgr2z4;
assign vis_psp_o[10] = Oir2z4;
assign Cfdvx4 = Dkr2z4;
assign Ngdvx4 = Slr2z4;
assign vis_r1_o[13] = Hnr2z4;
assign vis_r5_o[13] = Wor2z4;
assign vis_r7_o[13] = Lqr2z4;
assign vis_r1_o[8] = Asr2z4;
assign vis_r5_o[8] = Otr2z4;
assign vis_r7_o[8] = Cvr2z4;
assign vis_msp_o[6] = Qwr2z4;
assign vis_psp_o[6] = Eyr2z4;
assign M9dvx4 = Szr2z4;
assign Wadvx4 = G1s2z4;
assign vis_r1_o[9] = U2s2z4;
assign vis_r5_o[9] = I4s2z4;
assign vis_r7_o[9] = W5s2z4;
assign vis_r1_o[10] = K7s2z4;
assign vis_r5_o[10] = Z8s2z4;
assign vis_r7_o[10] = Oas2z4;
assign vis_msp_o[8] = Dcs2z4;
assign vis_psp_o[8] = Rds2z4;
assign Z7hvx4 = Ffs2z4;
assign Zuh2z4[27] = Vgs2z4;
assign Zuh2z4[26] = Mis2z4;
assign Zuh2z4[28] = Dks2z4;
assign Zuh2z4[29] = Uls2z4;
assign Zuh2z4[30] = Lns2z4;
assign Zuh2z4[31] = Cps2z4;
assign Zuh2z4[19] = Tqs2z4;
assign Zuh2z4[18] = Kss2z4;
assign Zuh2z4[20] = Bus2z4;
assign Zuh2z4[21] = Svs2z4;
assign Zuh2z4[22] = Jxs2z4;
assign Zuh2z4[23] = Azs2z4;
assign Eg8vx4 = R0t2z4;
assign Ot9vx4 = I2t2z4;
assign Dmgvx4 = A4t2z4;
assign Fjgvx4 = O5t2z4;
assign Q5gvx4 = Y6t2z4;
assign Mj8vx4 = L8t2z4;
assign Pp8vx4 = Y9t2z4;
assign Nngvx4 = Mbt2z4;
assign Vogvx4 = Adt2z4;
assign Hx8vx4 = Pet2z4;
assign vis_r6_o[31] = Cgt2z4;
assign vis_r6_o[28] = Rht2z4;
assign vis_r6_o[7] = Gjt2z4;
assign vis_r6_o[1] = Ukt2z4;
assign vis_r6_o[0] = Imt2z4;
assign vis_r6_o[30] = Wnt2z4;
assign vis_r6_o[29] = Lpt2z4;
assign vis_r6_o[27] = Art2z4;
assign vis_r6_o[26] = Pst2z4;
assign vis_r6_o[25] = Eut2z4;
assign vis_r6_o[24] = Tvt2z4;
assign vis_r6_o[6] = Ixt2z4;
assign vis_r6_o[5] = Wyt2z4;
assign vis_r6_o[4] = K0u2z4;
assign vis_r6_o[3] = Y1u2z4;
assign vis_r6_o[22] = M3u2z4;
assign vis_r6_o[21] = B5u2z4;
assign vis_r6_o[19] = Q6u2z4;
assign vis_r6_o[18] = F8u2z4;
assign vis_r6_o[17] = U9u2z4;
assign vis_r6_o[16] = Jbu2z4;
assign vis_r6_o[14] = Ycu2z4;
assign vis_r6_o[13] = Neu2z4;
assign vis_r6_o[12] = Cgu2z4;
assign vis_r6_o[10] = Rhu2z4;
assign vis_r6_o[2] = Gju2z4;
assign vis_r6_o[9] = Uku2z4;
assign vis_r6_o[8] = Imu2z4;
assign vis_r6_o[15] = Wnu2z4;
assign vis_r4_o[31] = Lpu2z4;
assign vis_r4_o[28] = Aru2z4;
assign vis_r4_o[7] = Psu2z4;
assign vis_r4_o[1] = Duu2z4;
assign vis_r4_o[0] = Rvu2z4;
assign vis_r4_o[30] = Fxu2z4;
assign vis_r4_o[29] = Uyu2z4;
assign vis_r4_o[27] = J0v2z4;
assign vis_r4_o[26] = Y1v2z4;
assign vis_r4_o[25] = N3v2z4;
assign vis_r4_o[24] = C5v2z4;
assign vis_r4_o[6] = R6v2z4;
assign vis_r4_o[5] = F8v2z4;
assign vis_r4_o[4] = T9v2z4;
assign vis_r4_o[3] = Hbv2z4;
assign vis_r4_o[22] = Vcv2z4;
assign vis_r4_o[21] = Kev2z4;
assign vis_r4_o[19] = Zfv2z4;
assign vis_r4_o[18] = Ohv2z4;
assign vis_r4_o[17] = Djv2z4;
assign vis_r4_o[16] = Skv2z4;
assign vis_r4_o[14] = Hmv2z4;
assign vis_r4_o[13] = Wnv2z4;
assign vis_r4_o[12] = Lpv2z4;
assign vis_r4_o[10] = Arv2z4;
assign vis_r4_o[2] = Psv2z4;
assign vis_r4_o[9] = Duv2z4;
assign vis_r4_o[8] = Rvv2z4;
assign vis_r4_o[15] = Fxv2z4;
assign Wtgvx4 = Uyv2z4;
assign vis_ipsr_o[1] = G0w2z4;
assign vis_ipsr_o[0] = R1w2z4;
assign Zph2z4[0] = C3w2z4;
assign Rkgvx4 = S4w2z4;
assign Ul8vx4 = I6w2z4;
assign Krgvx4 = U7w2z4;
assign Ki8vx4 = G9w2z4;
assign Xyfvx4 = Vaw2z4;
assign Mxfvx4 = Jcw2z4;
assign Cbfvx4 = Ydw2z4;
assign Mcfvx4 = Mfw2z4;
assign Wdfvx4 = Ahw2z4;
assign Gffvx4 = Oiw2z4;
assign Qgfvx4 = Ckw2z4;
assign Aifvx4 = Qlw2z4;
assign Kjfvx4 = Enw2z4;
assign Ukfvx4 = Sow2z4;
assign Emfvx4 = Gqw2z4;
assign Onfvx4 = Urw2z4;
assign Yofvx4 = Itw2z4;
assign Jqfvx4 = Xuw2z4;
assign Urfvx4 = Mww2z4;
assign Ftfvx4 = Byw2z4;
assign Qufvx4 = Qzw2z4;
assign Bwfvx4 = F1x2z4;
assign Aj9vx4 = U2x2z4;
assign vis_pc_o[1] = J4x2z4;
assign Mk8vx4 = U5x2z4;
assign vis_pc_o[2] = G7x2z4;
assign vis_pc_o[3] = R8x2z4;
assign vis_pc_o[4] = Cax2z4;
assign vis_pc_o[5] = Nbx2z4;
assign vis_pc_o[6] = Ycx2z4;
assign vis_pc_o[7] = Jex2z4;
assign vis_pc_o[9] = Ufx2z4;
assign vis_pc_o[11] = Fhx2z4;
assign vis_pc_o[13] = Rix2z4;
assign vis_pc_o[15] = Dkx2z4;
assign vis_pc_o[16] = Plx2z4;
assign vis_pc_o[17] = Bnx2z4;
assign vis_pc_o[21] = Nox2z4;
assign vis_pc_o[24] = Zpx2z4;
assign vis_pc_o[25] = Lrx2z4;
assign vis_pc_o[26] = Xsx2z4;
assign vis_pc_o[27] = Jux2z4;
assign vis_pc_o[28] = Vvx2z4;
assign A3gvx4 = Hxx2z4;
assign I4gvx4 = Tyx2z4;
assign Fuevx4 = F0y2z4;
assign R9fvx4 = T1y2z4;
assign Pvevx4 = I3y2z4;
assign Zwevx4 = W4y2z4;
assign Jyevx4 = K6y2z4;
assign Tzevx4 = Y7y2z4;
assign D1fvx4 = M9y2z4;
assign O2fvx4 = Bby2z4;
assign Z3fvx4 = Qcy2z4;
assign V6fvx4 = Fey2z4;
assign G8fvx4 = Ufy2z4;
assign V8evx4 = Jhy2z4;
assign I29vx4 = Viy2z4;
assign P39vx4 = Jky2z4;
assign W49vx4 = Xly2z4;
assign D69vx4 = Lny2z4;
assign K79vx4 = Zoy2z4;
assign R89vx4 = Nqy2z4;
assign Y99vx4 = Bsy2z4;
assign Fb9vx4 = Pty2z4;
assign Mc9vx4 = Dvy2z4;
assign Ud9vx4 = Swy2z4;
assign Cf9vx4 = Hyy2z4;
assign Tjh2z4[2] = Wzy2z4;
assign Wv9vx4 = K1z2z4;
assign Bx9vx4 = C3z2z4;
assign Uzcvx4 = U4z2z4;
assign Cq9vx4 = I6z2z4;
assign Gr9vx4 = W7z2z4;
assign Ks9vx4 = K9z2z4;
assign Nt8vx4 = Yaz2z4;
assign vis_psp_o[5] = Mcz2z4;
assign vis_psp_o[26] = Aez2z4;
assign vis_psp_o[29] = Pfz2z4;
assign vis_r12_o[31] = Ehz2z4;
assign vis_r12_o[28] = Tiz2z4;
assign vis_r12_o[7] = Ikz2z4;
assign vis_r12_o[1] = Wlz2z4;
assign vis_r12_o[0] = Knz2z4;
assign vis_r12_o[29] = Yoz2z4;
assign vis_r12_o[26] = Nqz2z4;
assign vis_r12_o[25] = Csz2z4;
assign vis_r12_o[6] = Rtz2z4;
assign vis_r12_o[5] = Fvz2z4;
assign vis_r12_o[4] = Twz2z4;
assign vis_r12_o[3] = Hyz2z4;
assign vis_r12_o[22] = Vzz2z4;
assign vis_r12_o[18] = K103z4;
assign vis_r12_o[17] = Z203z4;
assign vis_r12_o[16] = O403z4;
assign vis_r12_o[14] = D603z4;
assign vis_r12_o[12] = S703z4;
assign vis_r12_o[10] = H903z4;
assign vis_r12_o[2] = Wa03z4;
assign vis_r12_o[8] = Kc03z4;
assign vis_r14_o[31] = Yd03z4;
assign vis_r14_o[28] = Nf03z4;
assign vis_r14_o[7] = Ch03z4;
assign vis_r14_o[1] = Qi03z4;
assign vis_r14_o[0] = Ek03z4;
assign vis_r14_o[29] = Sl03z4;
assign vis_r14_o[26] = Hn03z4;
assign vis_r14_o[25] = Wo03z4;
assign vis_r14_o[6] = Lq03z4;
assign vis_r14_o[5] = Zr03z4;
assign vis_r14_o[4] = Nt03z4;
assign vis_r14_o[3] = Bv03z4;
assign vis_r14_o[22] = Pw03z4;
assign vis_r14_o[18] = Ey03z4;
assign vis_r14_o[17] = Tz03z4;
assign vis_r14_o[16] = I113z4;
assign vis_r14_o[14] = X213z4;
assign vis_r14_o[12] = M413z4;
assign vis_r14_o[10] = B613z4;
assign vis_r14_o[2] = Q713z4;
assign vis_r14_o[8] = E913z4;
assign vis_r11_o[31] = Sa13z4;
assign vis_r11_o[28] = Hc13z4;
assign vis_r11_o[7] = Wd13z4;
assign vis_r11_o[1] = Kf13z4;
assign vis_r11_o[0] = Yg13z4;
assign vis_r11_o[30] = Mi13z4;
assign vis_r11_o[29] = Bk13z4;
assign vis_r11_o[27] = Ql13z4;
assign vis_r11_o[26] = Fn13z4;
assign vis_r11_o[25] = Uo13z4;
assign vis_r11_o[24] = Jq13z4;
assign vis_r11_o[6] = Yr13z4;
assign vis_r11_o[5] = Mt13z4;
assign vis_r11_o[4] = Av13z4;
assign vis_r11_o[3] = Ow13z4;
assign vis_r11_o[22] = Cy13z4;
assign vis_r11_o[21] = Rz13z4;
assign vis_r11_o[19] = G123z4;
assign vis_r11_o[18] = V223z4;
assign vis_r11_o[17] = K423z4;
assign vis_r11_o[16] = Z523z4;
assign vis_r11_o[14] = O723z4;
assign vis_r11_o[13] = D923z4;
assign vis_r11_o[12] = Sa23z4;
assign vis_r11_o[10] = Hc23z4;
assign vis_r11_o[2] = Wd23z4;
assign vis_r11_o[9] = Kf23z4;
assign vis_r11_o[8] = Yg23z4;
assign vis_r11_o[15] = Mi23z4;
assign vis_r10_o[31] = Bk23z4;
assign vis_r10_o[28] = Ql23z4;
assign vis_r10_o[7] = Fn23z4;
assign vis_r10_o[1] = To23z4;
assign vis_r10_o[0] = Hq23z4;
assign vis_r10_o[30] = Vr23z4;
assign vis_r10_o[29] = Kt23z4;
assign vis_r10_o[27] = Zu23z4;
assign vis_r10_o[26] = Ow23z4;
assign vis_r10_o[25] = Dy23z4;
assign vis_r10_o[24] = Sz23z4;
assign vis_r10_o[6] = H133z4;
assign vis_r10_o[5] = V233z4;
assign vis_r10_o[4] = J433z4;
assign vis_r10_o[3] = X533z4;
assign vis_r10_o[22] = L733z4;
assign vis_r10_o[21] = A933z4;
assign vis_r10_o[19] = Pa33z4;
assign vis_r10_o[18] = Ec33z4;
assign vis_r10_o[17] = Td33z4;
assign vis_r10_o[16] = If33z4;
assign vis_r10_o[14] = Xg33z4;
assign vis_r10_o[13] = Mi33z4;
assign vis_r10_o[12] = Bk33z4;
assign vis_r10_o[10] = Ql33z4;
assign vis_r10_o[2] = Fn33z4;
assign vis_r10_o[9] = To33z4;
assign vis_r10_o[8] = Hq33z4;
assign vis_r10_o[15] = Vr33z4;
assign vis_r9_o[31] = Kt33z4;
assign vis_r9_o[28] = Zu33z4;
assign vis_r9_o[7] = Ow33z4;
assign vis_r9_o[1] = Cy33z4;
assign vis_r9_o[0] = Qz33z4;
assign vis_r9_o[30] = E143z4;
assign vis_r9_o[29] = T243z4;
assign vis_r9_o[27] = I443z4;
assign vis_r9_o[26] = X543z4;
assign vis_r9_o[25] = M743z4;
assign vis_r9_o[24] = B943z4;
assign vis_r9_o[6] = Qa43z4;
assign vis_r9_o[5] = Ec43z4;
assign vis_r9_o[4] = Sd43z4;
assign vis_r9_o[3] = Gf43z4;
assign vis_r9_o[22] = Ug43z4;
assign vis_r9_o[21] = Ji43z4;
assign vis_r9_o[19] = Yj43z4;
assign vis_r9_o[18] = Nl43z4;
assign vis_r9_o[17] = Cn43z4;
assign vis_r9_o[16] = Ro43z4;
assign vis_r9_o[14] = Gq43z4;
assign vis_r9_o[13] = Vr43z4;
assign vis_r9_o[12] = Kt43z4;
assign vis_r9_o[10] = Zu43z4;
assign vis_r9_o[2] = Ow43z4;
assign vis_r9_o[9] = Cy43z4;
assign vis_r9_o[8] = Qz43z4;
assign vis_r9_o[15] = E153z4;
assign vis_r8_o[31] = T253z4;
assign vis_r8_o[28] = I453z4;
assign vis_r8_o[7] = X553z4;
assign vis_r8_o[1] = L753z4;
assign vis_r8_o[0] = Z853z4;
assign vis_r8_o[30] = Na53z4;
assign vis_r8_o[29] = Cc53z4;
assign vis_r8_o[27] = Rd53z4;
assign vis_r8_o[26] = Gf53z4;
assign vis_r8_o[25] = Vg53z4;
assign vis_r8_o[24] = Ki53z4;
assign vis_r8_o[6] = Zj53z4;
assign vis_r8_o[5] = Nl53z4;
assign vis_r8_o[4] = Bn53z4;
assign vis_r8_o[3] = Po53z4;
assign vis_r8_o[22] = Dq53z4;
assign vis_r8_o[21] = Sr53z4;
assign vis_r8_o[19] = Ht53z4;
assign vis_r8_o[18] = Wu53z4;
assign vis_r8_o[17] = Lw53z4;
assign vis_r8_o[16] = Ay53z4;
assign vis_r8_o[14] = Pz53z4;
assign vis_r8_o[13] = E163z4;
assign vis_r8_o[12] = T263z4;
assign vis_r8_o[10] = I463z4;
assign vis_r8_o[2] = X563z4;
assign vis_r8_o[9] = L763z4;
assign vis_r8_o[8] = Z863z4;
assign vis_r8_o[15] = Na63z4;
assign vis_r3_o[31] = Cc63z4;
assign vis_r3_o[28] = Rd63z4;
assign vis_r3_o[7] = Gf63z4;
assign vis_r3_o[1] = Ug63z4;
assign vis_r3_o[0] = Ii63z4;
assign vis_r3_o[30] = Wj63z4;
assign vis_r3_o[29] = Ll63z4;
assign vis_r3_o[27] = An63z4;
assign vis_r3_o[26] = Po63z4;
assign vis_r3_o[25] = Eq63z4;
assign vis_r3_o[24] = Tr63z4;
assign vis_r3_o[6] = It63z4;
assign vis_r3_o[5] = Wu63z4;
assign vis_r3_o[4] = Kw63z4;
assign vis_r3_o[3] = Yx63z4;
assign vis_r3_o[22] = Mz63z4;
assign vis_r3_o[21] = B173z4;
assign vis_r3_o[19] = Q273z4;
assign vis_r3_o[18] = F473z4;
assign vis_r3_o[17] = U573z4;
assign vis_r3_o[16] = J773z4;
assign vis_r3_o[14] = Y873z4;
assign vis_r3_o[13] = Na73z4;
assign vis_r3_o[12] = Cc73z4;
assign vis_r3_o[10] = Rd73z4;
assign vis_r3_o[2] = Gf73z4;
assign vis_r3_o[9] = Ug73z4;
assign vis_r3_o[8] = Ii73z4;
assign vis_r3_o[15] = Wj73z4;
assign vis_r2_o[31] = Ll73z4;
assign vis_r2_o[28] = An73z4;
assign vis_r2_o[7] = Po73z4;
assign vis_r2_o[1] = Dq73z4;
assign vis_r2_o[0] = Rr73z4;
assign vis_r2_o[30] = Ft73z4;
assign vis_r2_o[29] = Uu73z4;
assign vis_r2_o[27] = Jw73z4;
assign vis_r2_o[26] = Yx73z4;
assign vis_r2_o[25] = Nz73z4;
assign vis_r2_o[24] = C183z4;
assign vis_r2_o[6] = R283z4;
assign vis_r2_o[5] = F483z4;
assign vis_r2_o[4] = T583z4;
assign vis_r2_o[3] = H783z4;
assign vis_r2_o[22] = V883z4;
assign vis_r2_o[21] = Ka83z4;
assign vis_r2_o[19] = Zb83z4;
assign vis_r2_o[18] = Od83z4;
assign vis_r2_o[17] = Df83z4;
assign vis_r2_o[16] = Sg83z4;
assign vis_r2_o[14] = Hi83z4;
assign vis_r2_o[13] = Wj83z4;
assign vis_r2_o[12] = Ll83z4;
assign vis_r2_o[10] = An83z4;
assign vis_r2_o[2] = Po83z4;
assign vis_r2_o[9] = Dq83z4;
assign vis_r2_o[8] = Rr83z4;
assign vis_r2_o[15] = Ft83z4;
assign vis_r0_o[30] = Uu83z4;
assign vis_r0_o[29] = Jw83z4;
assign vis_r0_o[27] = Yx83z4;
assign vis_r0_o[26] = Nz83z4;
assign vis_r0_o[25] = C193z4;
assign vis_r0_o[24] = R293z4;
assign vis_r0_o[6] = G493z4;
assign S6dvx4 = U593z4;
assign C8dvx4 = I793z4;
assign vis_r0_o[5] = W893z4;
assign vis_r0_o[4] = Ka93z4;
assign vis_r0_o[3] = Yb93z4;
assign vis_r0_o[22] = Md93z4;
assign vis_r0_o[21] = Bf93z4;
assign vis_r0_o[19] = Qg93z4;
assign vis_r0_o[18] = Fi93z4;
assign vis_r0_o[17] = Uj93z4;
assign vis_r0_o[16] = Jl93z4;
assign Ukdvx4 = Ym93z4;
assign vis_r0_o[14] = No93z4;
assign vis_r0_o[13] = Cq93z4;
assign vis_r0_o[12] = Rr93z4;
assign vis_r0_o[10] = Gt93z4;
assign vis_r0_o[2] = Vu93z4;
assign E1dvx4 = Jw93z4;
assign O2dvx4 = Xx93z4;
assign N6hvx4 = Lz93z4;
assign Uth2z4[0] = B1a3z4;
assign Uth2z4[1] = P2a3z4;
assign Czh2z4[15] = D4a3z4;
assign Czh2z4[14] = U5a3z4;
assign Czh2z4[12] = L7a3z4;
assign Czh2z4[10] = C9a3z4;
assign Czh2z4[4] = Taa3z4;
assign Czh2z4[23] = Jca3z4;
assign Czh2z4[0] = Aea3z4;
assign Czh2z4[1] = Qfa3z4;
assign Czh2z4[2] = Gha3z4;
assign Czh2z4[3] = Wia3z4;
assign Czh2z4[5] = Mka3z4;
assign Czh2z4[22] = Cma3z4;
assign F2hvx4 = Tna3z4;
assign Irh2z4[19] = Jpa3z4;
assign Irh2z4[15] = Ara3z4;
assign Irh2z4[14] = Rsa3z4;
assign Irh2z4[12] = Iua3z4;
assign Irh2z4[10] = Zva3z4;
assign Irh2z4[5] = Qxa3z4;
assign Irh2z4[4] = Gza3z4;
assign Irh2z4[3] = W0b3z4;
assign Irh2z4[2] = M2b3z4;
assign Irh2z4[1] = C4b3z4;
assign S0hvx4 = S5b3z4;
assign Czh2z4[6] = J7b3z4;
assign Irh2z4[6] = Z8b3z4;
assign Zuh2z4[24] = Pab3z4;
assign Zuh2z4[16] = Gcb3z4;
assign Zuh2z4[8] = Xdb3z4;
assign Czh2z4[7] = Nfb3z4;
assign Irh2z4[7] = Dhb3z4;
assign Zuh2z4[25] = Tib3z4;
assign Zuh2z4[17] = Kkb3z4;
assign Zuh2z4[9] = Bmb3z4;
assign D3i2z4[4] = Rnb3z4;
assign T1i2z4[4] = Ipb3z4;
assign D3i2z4[0] = Zqb3z4;
assign D3i2z4[3] = Qsb3z4;
assign T1i2z4[3] = Hub3z4;
assign D3i2z4[2] = Yvb3z4;
assign T1i2z4[2] = Pxb3z4;
assign D3i2z4[7] = Gzb3z4;
assign T1i2z4[7] = X0c3z4;
assign D3i2z4[6] = O2c3z4;
assign T1i2z4[6] = F4c3z4;
assign D3i2z4[5] = W5c3z4;
assign T1i2z4[5] = N7c3z4;
assign D3i2z4[1] = E9c3z4;
assign T1i2z4[1] = Vac3z4;
assign L0i2z4[1] = Mcc3z4;
assign L0i2z4[2] = Bec3z4;
assign L0i2z4[3] = Qfc3z4;
assign L0i2z4[4] = Fhc3z4;
assign L0i2z4[5] = Uic3z4;
assign L0i2z4[6] = Jkc3z4;
assign L0i2z4[7] = Ylc3z4;
assign L0i2z4[10] = Nnc3z4;
assign L0i2z4[12] = Dpc3z4;
assign L0i2z4[14] = Tqc3z4;
assign L0i2z4[15] = Jsc3z4;
assign L0i2z4[0] = Ztc3z4;
assign Y3dvx4 = Ovc3z4;
assign vis_r0_o[9] = Cxc3z4;
assign vis_r0_o[8] = Qyc3z4;
assign vis_r0_o[15] = E0d3z4;
assign Vu8vx4 = T1d3z4;
assign Fs8vx4 = H3d3z4;
assign vis_pc_o[8] = V4d3z4;
assign Oy8vx4 = G6d3z4;
assign Zuh2z4[3] = T7d3z4;
assign Zuh2z4[0] = J9d3z4;
assign Zuh2z4[1] = Zad3z4;
assign Zuh2z4[2] = Pcd3z4;
assign Zuh2z4[4] = Fed3z4;
assign Zuh2z4[5] = Vfd3z4;
assign Zuh2z4[6] = Lhd3z4;
assign Zuh2z4[7] = Bjd3z4;
assign Gcdvx4 = Rkd3z4;
assign vis_pc_o[10] = Gmd3z4;
assign vis_r0_o[11] = Snd3z4;
assign vis_r1_o[11] = Hpd3z4;
assign vis_r2_o[11] = Wqd3z4;
assign vis_r3_o[11] = Lsd3z4;
assign vis_r8_o[11] = Aud3z4;
assign vis_r9_o[11] = Pvd3z4;
assign vis_r10_o[11] = Exd3z4;
assign vis_r11_o[11] = Tyd3z4;
assign vis_r4_o[11] = I0e3z4;
assign vis_r5_o[11] = X1e3z4;
assign vis_r6_o[11] = M3e3z4;
assign vis_r7_o[11] = B5e3z4;
assign vis_r12_o[11] = Q6e3z4;
assign vis_r14_o[11] = F8e3z4;
assign vis_msp_o[9] = U9e3z4;
assign vis_psp_o[9] = Ibe3z4;
assign Rddvx4 = Wce3z4;
assign L0i2z4[11] = Lee3z4;
assign Czh2z4[11] = Bge3z4;
assign Irh2z4[11] = She3z4;
assign D3i2z4[11] = Jje3z4;
assign T1i2z4[11] = Ble3z4;
assign vis_pc_o[12] = Tme3z4;
assign vis_pc_o[20] = Foe3z4;
assign vis_r12_o[9] = Rpe3z4;
assign vis_r14_o[9] = Fre3z4;
assign vis_msp_o[7] = Tse3z4;
assign vis_psp_o[7] = Hue3z4;
assign L0i2z4[9] = Vve3z4;
assign Czh2z4[9] = Kxe3z4;
assign Irh2z4[9] = Aze3z4;
assign D3i2z4[9] = Q0f3z4;
assign L0i2z4[8] = H2f3z4;
assign Czh2z4[8] = W3f3z4;
assign Irh2z4[8] = M5f3z4;
assign D3i2z4[8] = C7f3z4;
assign T1i2z4[8] = T8f3z4;
assign vis_pc_o[22] = Kaf3z4;
assign vis_r0_o[23] = Wbf3z4;
assign vis_r2_o[23] = Ldf3z4;
assign vis_r3_o[23] = Aff3z4;
assign vis_r8_o[23] = Pgf3z4;
assign vis_r9_o[23] = Eif3z4;
assign vis_r10_o[23] = Tjf3z4;
assign vis_r11_o[23] = Ilf3z4;
assign vis_r4_o[23] = Xmf3z4;
assign vis_r5_o[23] = Mof3z4;
assign vis_r6_o[23] = Bqf3z4;
assign vis_r12_o[23] = Qrf3z4;
assign vis_r14_o[23] = Ftf3z4;
assign vis_psp_o[21] = Uuf3z4;
assign vis_pc_o[14] = Jwf3z4;
assign vis_r12_o[13] = Vxf3z4;
assign vis_r14_o[13] = Kzf3z4;
assign vis_msp_o[11] = Z0g3z4;
assign vis_psp_o[11] = O2g3z4;
assign L0i2z4[13] = D4g3z4;
assign Czh2z4[13] = T5g3z4;
assign Irh2z4[13] = K7g3z4;
assign vis_pc_o[19] = B9g3z4;
assign vis_r0_o[20] = Nag3z4;
assign vis_r1_o[20] = Ccg3z4;
assign vis_r2_o[20] = Rdg3z4;
assign vis_r3_o[20] = Gfg3z4;
assign vis_r8_o[20] = Vgg3z4;
assign vis_r9_o[20] = Kig3z4;
assign vis_r10_o[20] = Zjg3z4;
assign vis_r11_o[20] = Olg3z4;
assign vis_r4_o[20] = Dng3z4;
assign vis_r5_o[20] = Sog3z4;
assign vis_r6_o[20] = Hqg3z4;
assign vis_r7_o[20] = Wrg3z4;
assign vis_r12_o[20] = Ltg3z4;
assign vis_r14_o[20] = Avg3z4;
assign vis_msp_o[18] = Pwg3z4;
assign vis_psp_o[18] = Eyg3z4;
assign Mqdvx4 = Tzg3z4;
assign Czh2z4[20] = I1h3z4;
assign Irh2z4[20] = Z2h3z4;
assign D3i2z4[14] = Q4h3z4;
assign D3i2z4[15] = I6h3z4;
assign vis_r12_o[21] = A8h3z4;
assign vis_r14_o[21] = P9h3z4;
assign vis_msp_o[19] = Ebh3z4;
assign vis_psp_o[19] = Tch3z4;
assign Czh2z4[21] = Ieh3z4;
assign Itdvx4 = Zfh3z4;
assign W1evx4 = Ohh3z4;
assign vis_r12_o[27] = Djh3z4;
assign vis_r14_o[27] = Skh3z4;
assign vis_msp_o[25] = Hmh3z4;
assign vis_psp_o[25] = Wnh3z4;
assign vis_r12_o[15] = Lph3z4;
assign vis_r14_o[15] = Arh3z4;
assign vis_msp_o[13] = Psh3z4;
assign vis_psp_o[13] = Euh3z4;
assign vis_r12_o[19] = Tvh3z4;
assign vis_r14_o[19] = Ixh3z4;
assign vis_msp_o[17] = Xyh3z4;
assign vis_psp_o[17] = M0i3z4;
assign Czh2z4[17] = B2i3z4;
assign Irh2z4[17] = S3i3z4;
assign vis_r12_o[30] = J5i3z4;
assign vis_r14_o[30] = Y6i3z4;
assign vis_msp_o[28] = N8i3z4;
assign vis_psp_o[28] = Cai3z4;
assign H0gvx4 = Rbi3z4;
assign Irh2z4[22] = Ddi3z4;
assign Irh2z4[23] = Uei3z4;
assign Pxdvx4 = Lgi3z4;
assign Cvgvx4 = Aii3z4;
assign vis_r12_o[24] = Qji3z4;
assign vis_r14_o[24] = Fli3z4;
assign vis_msp_o[22] = Umi3z4;
assign vis_psp_o[22] = Joi3z4;
assign sys_reset_req_o = Ypi3z4;
assign Jchvx4 = (!Ypi3z4);
assign Iwh2z4 = (Irh2z4 - 1'b1);
assign {Enh2z4, N4i2z4} = ({Lkevx4, Zievx4, Nhevx4, Bgevx4, Peevx4, 
 Ddevx4, Rbevx4, Faevx4, A3ivx4} - 1'b1);
assign Roh2z4 = (vis_pc_o + 1'b1);
assign {Ykh2z4, L5i2z4} = ({vis_pc_o[30:2], P1gvx4} + 1'b1);
assign Pri3z4 = ({{Jz9vx4, M0avx4, P1avx4, S2avx4, V3avx4, Y4avx4,
 B6avx4, E7avx4, H8avx4, K9avx4, Naavx4, Qbavx4, Tcavx4, Wdavx4,
 Zeavx4, Cgavx4, Fhavx4, Iiavx4, Ljavx4, Okavx4, Rlavx4, Umavx4,
 Xnavx4, Apavx4, Dqavx4, Gravx4, Jsavx4, Ltavx4, Nuavx4, Pvavx4,
 Rwavx4, Txavx4, Vyavx4}, 1'b0} + {{1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Xzavx4}, 1'b1});
assign {Gy9vx4, Dmh2z4} = Pri3z4[33:1];
assign Fti3z4 = ({{1'b0, Zwcvx4, Ovcvx4, Ducvx4, Sscvx4, Hrcvx4, Wpcvx4,
 Locvx4, Ancvx4, Plcvx4, Ekcvx4, Ticvx4, Ihcvx4, Xfcvx4, Mecvx4,
 Bdcvx4, Qbcvx4, Facvx4, U8cvx4, J7cvx4, Y5cvx4, N4cvx4, C3cvx4,
 S1cvx4, I0cvx4, Yybvx4, Oxbvx4, Ewbvx4, Uubvx4, Ktbvx4, Asbvx4,
 Qqbvx4, Gpbvx4}, 1'b0} + {{1'b0, Phh2z4, Dih2z4, Kih2z4, Whh2z4,
 Yih2z4, Vnbvx4, Kmbvx4, Rih2z4, Fjh2z4, Zkbvx4, Ojbvx4, Dibvx4,
 Sgbvx4, Hfbvx4, Wdbvx4, Lcbvx4, Abbvx4, P9bvx4, E8bvx4, T6bvx4,
 I5bvx4, Mjh2z4, Bhh2z4, Y3bvx4, Ugh2z4, O2bvx4, Zfh2z4, Ggh2z4,
 Sfh2z4, Ngh2z4, Ihh2z4, E1bvx4}, 1'b1});
assign {Jz9vx4, M0avx4, P1avx4, S2avx4, V3avx4, Y4avx4, B6avx4, E7avx4, 
 H8avx4, K9avx4, Naavx4, Qbavx4, Tcavx4, Wdavx4, Zeavx4, Cgavx4, 
 Fhavx4, Iiavx4, Ljavx4, Okavx4, Rlavx4, Umavx4, Xnavx4, Apavx4, 
 Dqavx4, Gravx4, Jsavx4, Ltavx4, Nuavx4, Pvavx4, Rwavx4, Txavx4, 
 Vyavx4} = Fti3z4[33:1];
assign Lkevx4 = (K5fvx4 & Xlevx4);
assign Zievx4 = (Z3fvx4 & Xlevx4);
assign Nhevx4 = (O2fvx4 & Xlevx4);
assign Bgevx4 = (D1fvx4 & Xlevx4);
assign Peevx4 = (Tzevx4 & Xlevx4);
assign Ddevx4 = (Jyevx4 & Xlevx4);
assign Rbevx4 = (Zwevx4 & Xlevx4);
assign Faevx4 = (Pvevx4 & Xlevx4);
assign P1gvx4 = (~(Bnnvx4 & Innvx4));
assign Innvx4 = (Pnnvx4 | Wnnvx4);
assign S1cvx4 = (Donvx4 & Konvx4);
assign I0cvx4 = (Donvx4 & Ronvx4);
assign Yybvx4 = (Yonvx4 & Donvx4);
assign Oxbvx4 = (Donvx4 & Fpnvx4);
assign Ewbvx4 = (Mpnvx4 & Donvx4);
assign Uubvx4 = (Tpnvx4 & Donvx4);
assign Ktbvx4 = (Aqnvx4 & Donvx4);
assign Ovcvx4 = (Donvx4 & Hqnvx4);
assign Asbvx4 = (Oqnvx4 & Vqnvx4);
assign Vqnvx4 = (~(Crnvx4 & O8gvx4));
assign Crnvx4 = (~(Jrnvx4 | Mcgvx4));
assign Oqnvx4 = (Donvx4 & Qrnvx4);
assign Ducvx4 = (Xrnvx4 & Donvx4);
assign Sscvx4 = (Esnvx4 & Donvx4);
assign Hrcvx4 = (Lsnvx4 & Donvx4);
assign Wpcvx4 = (Donvx4 & Ssnvx4);
assign Locvx4 = (Donvx4 & Zsnvx4);
assign Ancvx4 = (Gtnvx4 & Donvx4);
assign Plcvx4 = (Ntnvx4 & Donvx4);
assign Ekcvx4 = (Donvx4 & Utnvx4);
assign Ticvx4 = (Donvx4 & Bunvx4);
assign Ihcvx4 = (Donvx4 & Iunvx4);
assign Qqbvx4 = (Punvx4 & Donvx4);
assign Xfcvx4 = (Donvx4 & Wunvx4);
assign Mecvx4 = (Donvx4 & Dvnvx4);
assign Bdcvx4 = (Donvx4 & Kvnvx4);
assign Qbcvx4 = (Donvx4 & Rvnvx4);
assign Facvx4 = (Donvx4 & Yvnvx4);
assign U8cvx4 = (Donvx4 & Fwnvx4);
assign J7cvx4 = (Donvx4 & Mwnvx4);
assign Y5cvx4 = (Donvx4 & Twnvx4);
assign N4cvx4 = (Donvx4 & Axnvx4);
assign C3cvx4 = (Hxnvx4 & Donvx4);
assign Gpbvx4 = (Donvx4 & Oxnvx4);
assign Xzavx4 = (O8gvx4 & Vxnvx4);
assign Vxnvx4 = (~(Cynvx4 & Jynvx4));
assign Jynvx4 = (Qynvx4 & Xynvx4);
assign Xynvx4 = (~(Eznvx4 & Lznvx4));
assign Lznvx4 = (~(Sznvx4 & Zznvx4));
assign Zznvx4 = (~(G0ovx4 & N0ovx4));
assign N0ovx4 = (~(U0ovx4 | B1ovx4));
assign Qynvx4 = (~(Cn8vx4 & I1ovx4));
assign I1ovx4 = (~(P1ovx4 & W1ovx4));
assign W1ovx4 = (~(D2ovx4 & U9gvx4));
assign P1ovx4 = (K2ovx4 | R2ovx4);
assign K2ovx4 = (M3ovx4 ? F3ovx4 : Y2ovx4);
assign Cynvx4 = (T3ovx4 & A4ovx4);
assign A4ovx4 = (H4ovx4 | Vdgvx4);
assign sleeping_o = (Cvgvx4 & O4ovx4);
assign Umnvx4 = (C5ovx4 ? V4ovx4 : Czh2z4[23]);
assign Nmnvx4 = (~(J5ovx4 & Q5ovx4));
assign Q5ovx4 = (X5ovx4 | hready_i);
assign J5ovx4 = (E6ovx4 & L6ovx4);
assign E6ovx4 = (~(S6ovx4 & Z6ovx4));
assign Gmnvx4 = (G7ovx4 & irq_i[0]);
assign G7ovx4 = (N7ovx4 & U7ovx4);
assign U7ovx4 = (~(B8ovx4 & I8ovx4));
assign N7ovx4 = (~(P8ovx4 & W8ovx4));
assign W8ovx4 = (D9ovx4 | K9ovx4);
assign P8ovx4 = (R9ovx4 & Y9ovx4);
assign R9ovx4 = (Faovx4 | hwdata_o[0]);
assign Faovx4 = (~(Maovx4 | Taovx4));
assign Zlnvx4 = (~(Abovx4 & Hbovx4));
assign Hbovx4 = (~(Xlevx4 & Obovx4));
assign Obovx4 = (Vbovx4 | Ccovx4);
assign Slnvx4 = (Jcovx4 | Qcovx4);
assign Jcovx4 = (Edovx4 ? R9fvx4 : Xcovx4);
assign Llnvx4 = (Ldovx4 | Sdovx4);
assign Sdovx4 = (Geovx4 ? Ho8vx4 : Zdovx4);
assign Zdovx4 = (~(Neovx4 | Ueovx4));
assign Ldovx4 = (~(Bfovx4 & Ifovx4));
assign Ifovx4 = (~(Mxfvx4 & Pfovx4));
assign Bfovx4 = (~(Wfovx4 & R9fvx4));
assign Elnvx4 = (~(Dgovx4 & Kgovx4));
assign Kgovx4 = (Rgovx4 | hready_i);
assign Dgovx4 = (Ygovx4 & L6ovx4);
assign Ygovx4 = (~(S6ovx4 & Fhovx4));
assign Fhovx4 = (haddr_o[7] | haddr_o[2]);
assign Xknvx4 = (~(Mhovx4 & Thovx4));
assign Thovx4 = (Aiovx4 | hready_i);
assign Mhovx4 = (Hiovx4 & L6ovx4);
assign Hiovx4 = (~(S6ovx4 & Oiovx4));
assign Oiovx4 = (haddr_o[5] | haddr_o[3]);
assign Qknvx4 = (~(Viovx4 & Cjovx4));
assign Cjovx4 = (Jjovx4 | hready_i);
assign Viovx4 = (Qjovx4 & L6ovx4);
assign Qjovx4 = (~(S6ovx4 & Xjovx4));
assign Xjovx4 = (~(Ekovx4 ^ haddr_o[10]));
assign Jknvx4 = (~(Lkovx4 & Skovx4));
assign Skovx4 = (Zkovx4 | hready_i);
assign Lkovx4 = (Glovx4 & L6ovx4);
assign L6ovx4 = (~(S6ovx4 & Nlovx4));
assign Nlovx4 = (~(Ulovx4 & Bmovx4));
assign Bmovx4 = (Imovx4 & Pmovx4);
assign Pmovx4 = (Wmovx4 & Dnovx4);
assign Dnovx4 = (Knovx4 & Rnovx4);
assign Knovx4 = (~(haddr_o[26] | haddr_o[27]));
assign Wmovx4 = (~(haddr_o[23] | haddr_o[24]));
assign Imovx4 = (Ynovx4 & Foovx4);
assign Foovx4 = (~(haddr_o[21] | haddr_o[22]));
assign Ynovx4 = (~(haddr_o[19] | haddr_o[20]));
assign Ulovx4 = (Moovx4 & Toovx4);
assign Toovx4 = (Apovx4 & Hpovx4);
assign Hpovx4 = (Opovx4 & Vpovx4);
assign Opovx4 = (~(haddr_o[17] | haddr_o[18]));
assign Apovx4 = (haddr_o[15] & Cqovx4);
assign Moovx4 = (Jqovx4 & Qqovx4);
assign Qqovx4 = (haddr_o[14] & hsize_o[1]);
assign Jqovx4 = (Xqovx4 & haddr_o[13]);
assign Xqovx4 = (~(Erovx4 & Lrovx4));
assign Lrovx4 = (~(Srovx4 & Zrovx4));
assign Zrovx4 = (Gsovx4 & Ekovx4);
assign Gsovx4 = (Nsovx4 | Usovx4);
assign Srovx4 = (Btovx4 & Itovx4);
assign Itovx4 = (haddr_o[8] ^ haddr_o[9]);
assign Btovx4 = (haddr_o[11] ? Wtovx4 : Ptovx4);
assign Wtovx4 = (Duovx4 & haddr_o[10]);
assign Ptovx4 = (Kuovx4 & Nsovx4);
assign Nsovx4 = (Ruovx4 & Yuovx4);
assign Ruovx4 = (~(haddr_o[6] | haddr_o[2]));
assign haddr_o[2] = (!Fvovx4);
assign Kuovx4 = (~(haddr_o[10] | haddr_o[5]));
assign Erovx4 = (Mvovx4 | Tvovx4);
assign Tvovx4 = (haddr_o[8] ? Awovx4 : haddr_o[11]);
assign haddr_o[8] = (!Z6ovx4);
assign Awovx4 = (~(Hwovx4 & haddr_o[10]));
assign Hwovx4 = (~(Fvovx4 | Owovx4));
assign haddr_o[11] = (!Owovx4);
assign Mvovx4 = (~(Usovx4 & Vwovx4));
assign Vwovx4 = (~(Cxovx4 & Jxovx4));
assign Cxovx4 = (~(haddr_o[4] | haddr_o[3]));
assign haddr_o[3] = (!Ekovx4);
assign Usovx4 = (Qxovx4 & Duovx4);
assign Duovx4 = (~(haddr_o[7] | haddr_o[9]));
assign haddr_o[9] = (!Xxovx4);
assign Qxovx4 = (~(haddr_o[5] | haddr_o[6]));
assign Glovx4 = (~(S6ovx4 & Yuovx4));
assign Cknvx4 = (~(Eyovx4 & Lyovx4));
assign Lyovx4 = (~(L0i2z4[0] & Syovx4));
assign Syovx4 = (~(hwdata_o[0] & Zyovx4));
assign Eyovx4 = (~(Gzovx4 & hwdata_o[0]));
assign Vjnvx4 = (~(Nzovx4 & Uzovx4));
assign Uzovx4 = (B0pvx4 & I0pvx4);
assign I0pvx4 = (~(P0pvx4 & vis_tbit_o));
assign B0pvx4 = (~(vis_pc_o[23] & W0pvx4));
assign Nzovx4 = (D1pvx4 & K1pvx4);
assign K1pvx4 = (R1pvx4 | Y1pvx4);
assign D1pvx4 = (~(Ewdvx4 & F2pvx4));
assign Ojnvx4 = (M2pvx4 | T2pvx4);
assign T2pvx4 = (A3pvx4 & H3pvx4);
assign A3pvx4 = (~(Ccovx4 | O3pvx4));
assign M2pvx4 = (C4pvx4 ? vis_tbit_o : V3pvx4);
assign C4pvx4 = (J4pvx4 & Q4pvx4);
assign Q4pvx4 = (X4pvx4 | Ccovx4);
assign J4pvx4 = (~(E5pvx4 & L5pvx4));
assign L5pvx4 = (S5pvx4 & Z5pvx4);
assign E5pvx4 = (G6pvx4 & N6pvx4);
assign N6pvx4 = (~(U6pvx4 & B7pvx4));
assign B7pvx4 = (~(I7pvx4 | P7pvx4));
assign U6pvx4 = (W7pvx4 & D8pvx4);
assign D8pvx4 = (F3ovx4 | B1ovx4);
assign W7pvx4 = (Mcgvx4 | Fjgvx4);
assign V3pvx4 = (~(K8pvx4 & R8pvx4));
assign R8pvx4 = (~(Y8pvx4 & F9pvx4));
assign K8pvx4 = (~(Dmh2z4[0] & M9pvx4));
assign Hjnvx4 = (~(T9pvx4 & Aapvx4));
assign Aapvx4 = (Hapvx4 & Oapvx4);
assign Oapvx4 = (~(Vapvx4 & hrdata_i[15]));
assign Hapvx4 = (Cbpvx4 & Jbpvx4);
assign Jbpvx4 = (~(Bwfvx4 & Pfovx4));
assign Cbpvx4 = (~(Qbpvx4 & hrdata_i[31]));
assign T9pvx4 = (Xbpvx4 & Ecpvx4);
assign Ecpvx4 = (~(G8fvx4 & Wfovx4));
assign Xbpvx4 = (Lcpvx4 | Scpvx4);
assign Ajnvx4 = (~(Zcpvx4 & Gdpvx4));
assign Gdpvx4 = (Ndpvx4 & Udpvx4);
assign Udpvx4 = (~(hrdata_i[13] & Vapvx4));
assign Ndpvx4 = (Bepvx4 & Iepvx4);
assign Iepvx4 = (~(Ftfvx4 & Pfovx4));
assign Bepvx4 = (~(hrdata_i[29] & Qbpvx4));
assign Zcpvx4 = (Pepvx4 & Wepvx4);
assign Wepvx4 = (~(Wfovx4 & K5fvx4));
assign Pepvx4 = (Dfpvx4 | Scpvx4);
assign Tinvx4 = (Rfpvx4 ? Kfpvx4 : Ik9vx4);
assign Kfpvx4 = (~(Yfpvx4 & Fgpvx4));
assign Fgpvx4 = (Mgpvx4 & Tgpvx4);
assign Tgpvx4 = (Ahpvx4 & Hhpvx4);
assign Ahpvx4 = (~(Ohpvx4 | Vhpvx4));
assign Mgpvx4 = (Cipvx4 & Jipvx4);
assign Jipvx4 = (~(Qipvx4 & Xipvx4));
assign Qipvx4 = (Ejpvx4 ^ Ljpvx4);
assign Cipvx4 = (Sjpvx4 & Zjpvx4);
assign Zjpvx4 = (~(Gkpvx4 & Nkpvx4));
assign Gkpvx4 = (Ukpvx4 & Dfpvx4);
assign Sjpvx4 = (~(Blpvx4 & Ilpvx4));
assign Blpvx4 = (~(B1ovx4 | Nggvx4));
assign Yfpvx4 = (Plpvx4 & Wlpvx4);
assign Wlpvx4 = (Dmpvx4 & Kmpvx4);
assign Kmpvx4 = (~(Uz8vx4 & Rmpvx4));
assign Dmpvx4 = (Ympvx4 & Fnpvx4);
assign Fnpvx4 = (~(K79vx4 & Mnpvx4));
assign Ympvx4 = (Tnpvx4 | Aopvx4);
assign Plpvx4 = (Hopvx4 & Oopvx4);
assign Oopvx4 = (~(Vopvx4 & Cppvx4));
assign Hopvx4 = (Jppvx4 | Efgvx4);
assign Minvx4 = (Xppvx4 ? Qppvx4 : vis_r0_o[1]);
assign Finvx4 = (Lqpvx4 ? Eqpvx4 : vis_apsr_o[1]);
assign Lqpvx4 = (Sqpvx4 & hready_i);
assign Sqpvx4 = (Zqpvx4 | Grpvx4);
assign Eqpvx4 = (~(Nrpvx4 & Urpvx4));
assign Urpvx4 = (X4pvx4 | Bspvx4);
assign Nrpvx4 = (Ispvx4 & Pspvx4);
assign Pspvx4 = (~(Wspvx4 & Dtpvx4));
assign Ispvx4 = (Ktpvx4 | Rtpvx4);
assign Yhnvx4 = (~(Ytpvx4 & Fupvx4));
assign Fupvx4 = (Mupvx4 & Tupvx4);
assign Tupvx4 = (~(P0pvx4 & vis_apsr_o[1]));
assign Mupvx4 = (~(W0pvx4 & vis_pc_o[28]));
assign Ytpvx4 = (Avpvx4 & Hvpvx4);
assign Hvpvx4 = (R1pvx4 | Ovpvx4);
assign Avpvx4 = (~(H3evx4 & F2pvx4));
assign Rhnvx4 = (~(Vvpvx4 & Cwpvx4));
assign Cwpvx4 = (~(Jwpvx4 & Wspvx4));
assign Vvpvx4 = (Ccovx4 ? Xwpvx4 : Qwpvx4);
assign Qwpvx4 = (~(Expvx4 & Lxpvx4));
assign Lxpvx4 = (~(Sxpvx4 & Wspvx4));
assign Sxpvx4 = (!Zxpvx4);
assign Expvx4 = (Grpvx4 ? Nypvx4 : Gypvx4);
assign Nypvx4 = (Uypvx4 & Bzpvx4);
assign Bzpvx4 = (~(Izpvx4 & Pzpvx4));
assign Pzpvx4 = (X4pvx4 | Wzpvx4);
assign Uypvx4 = (D0qvx4 | K0qvx4);
assign D0qvx4 = (!Wzpvx4);
assign Gypvx4 = (R0qvx4 & Y0qvx4);
assign Y0qvx4 = (~(Zwcvx4 & Dmh2z4[31]));
assign R0qvx4 = (Phh2z4 ? Zwcvx4 : Dmh2z4[31]);
assign Khnvx4 = (~(F1qvx4 & M1qvx4));
assign M1qvx4 = (T1qvx4 & A2qvx4);
assign A2qvx4 = (~(vis_apsr_o[0] & P0pvx4));
assign T1qvx4 = (~(W0pvx4 & vis_pc_o[27]));
assign F1qvx4 = (H2qvx4 & O2qvx4);
assign O2qvx4 = (R1pvx4 | V2qvx4);
assign H2qvx4 = (~(W1evx4 & F2pvx4));
assign Dhnvx4 = (Xppvx4 ? C3qvx4 : vis_r0_o[28]);
assign Wgnvx4 = (Xppvx4 ? J3qvx4 : vis_r0_o[31]);
assign Pgnvx4 = (~(Q3qvx4 & X3qvx4));
assign X3qvx4 = (~(C8dvx4 & F2pvx4));
assign Q3qvx4 = (E4qvx4 & L4qvx4);
assign L4qvx4 = (~(vis_pc_o[6] & W0pvx4));
assign E4qvx4 = (R1pvx4 | S4qvx4);
assign Ignvx4 = (Xppvx4 ? Z4qvx4 : vis_r0_o[7]);
assign Bgnvx4 = (Xppvx4 ? G5qvx4 : vis_r0_o[0]);
assign Ufnvx4 = (U5qvx4 ? N5qvx4 : Zph2z4[0]);
assign Nfnvx4 = (~(B6qvx4 & I6qvx4));
assign I6qvx4 = (~(P6qvx4 & W6qvx4));
assign P6qvx4 = (U5qvx4 & D7qvx4);
assign B6qvx4 = (~(K7qvx4 & Ccovx4));
assign K7qvx4 = (~(R7qvx4 & Y7qvx4));
assign Y7qvx4 = (~(hresp_i & F8qvx4));
assign F8qvx4 = (~(M8qvx4 & T8qvx4));
assign T8qvx4 = (A9qvx4 & H9qvx4);
assign H9qvx4 = (~(O9qvx4 & V9qvx4));
assign V9qvx4 = (~(Caqvx4 & Jaqvx4));
assign Jaqvx4 = (~(Qaqvx4 & Xaqvx4));
assign Xaqvx4 = (~(Ebqvx4 & Lbqvx4));
assign Ebqvx4 = (Sbqvx4 & Zbqvx4);
assign Zbqvx4 = (Gcqvx4 | Mcgvx4);
assign Sbqvx4 = (~(Ncqvx4 & Ucqvx4));
assign Caqvx4 = (Bdqvx4 | Dbgvx4);
assign A9qvx4 = (Idqvx4 & Pdqvx4);
assign Idqvx4 = (~(Wdqvx4 & Deqvx4));
assign Deqvx4 = (~(Keqvx4 & Reqvx4));
assign Reqvx4 = (~(Yeqvx4 & Ffqvx4));
assign Yeqvx4 = (~(U9gvx4 | Fjgvx4));
assign M8qvx4 = (Mfqvx4 & Tfqvx4);
assign Tfqvx4 = (Agqvx4 | Bdqvx4);
assign Mfqvx4 = (Hgqvx4 & Ogqvx4);
assign Ogqvx4 = (~(Whgvx4 & Vgqvx4));
assign Vgqvx4 = (~(Chqvx4 & Jhqvx4));
assign Jhqvx4 = (Qhqvx4 | Mcgvx4);
assign Chqvx4 = (~(Xhqvx4 & Eiqvx4));
assign Hgqvx4 = (~(P7pvx4 & Liqvx4));
assign Gfnvx4 = (Siqvx4 ? J3qvx4 : vis_r1_o[31]);
assign Zenvx4 = (Siqvx4 ? C3qvx4 : vis_r1_o[28]);
assign Senvx4 = (Siqvx4 ? Z4qvx4 : vis_r1_o[7]);
assign Lenvx4 = (Siqvx4 ? Qppvx4 : vis_r1_o[1]);
assign Eenvx4 = (Siqvx4 ? G5qvx4 : vis_r1_o[0]);
assign Xdnvx4 = (~(Ziqvx4 & Gjqvx4));
assign Ziqvx4 = (hready_i ? Ujqvx4 : Njqvx4);
assign Njqvx4 = (!vis_primask_o);
assign Qdnvx4 = (~(Bkqvx4 & Ikqvx4));
assign Ikqvx4 = (Pkqvx4 & Wkqvx4);
assign Wkqvx4 = (~(Vapvx4 & hrdata_i[0]));
assign Pkqvx4 = (Dlqvx4 & Klqvx4);
assign Klqvx4 = (~(Cbfvx4 & Pfovx4));
assign Dlqvx4 = (~(Qbpvx4 & hrdata_i[16]));
assign Bkqvx4 = (Rlqvx4 & Ylqvx4);
assign Ylqvx4 = (~(Hnevx4 & Wfovx4));
assign Rlqvx4 = (~(Uz8vx4 & Geovx4));
assign Jdnvx4 = (Rfpvx4 ? Fmqvx4 : Ml9vx4);
assign Fmqvx4 = (~(Mmqvx4 & Tmqvx4));
assign Tmqvx4 = (Anqvx4 & Hnqvx4);
assign Hnqvx4 = (Onqvx4 & Hhpvx4);
assign Onqvx4 = (~(Vnqvx4 & Xipvx4));
assign Vnqvx4 = (Coqvx4 ^ Joqvx4);
assign Anqvx4 = (Qoqvx4 & Xoqvx4);
assign Xoqvx4 = (~(Epqvx4 & Vopvx4));
assign Epqvx4 = (Lpqvx4 | Spqvx4);
assign Qoqvx4 = (~(Zpqvx4 & Uz8vx4));
assign Mmqvx4 = (Gqqvx4 & Nqqvx4);
assign Nqqvx4 = (Uqqvx4 & Brqvx4);
assign Brqvx4 = (~(Roevx4 & Irqvx4));
assign Uqqvx4 = (~(R89vx4 & Mnpvx4));
assign Gqqvx4 = (Prqvx4 & Wrqvx4);
assign Wrqvx4 = (~(B19vx4 & Rmpvx4));
assign Prqvx4 = (~(Dsqvx4 & K79vx4));
assign Cdnvx4 = (~(Ksqvx4 & Rsqvx4));
assign Rsqvx4 = (~(Ysqvx4 & Ftqvx4));
assign Ftqvx4 = (Mtqvx4 | Ttqvx4);
assign Ttqvx4 = (~(Auqvx4 | Huqvx4));
assign Ysqvx4 = (~(Ccovx4 | Abovx4));
assign Ksqvx4 = (O4ovx4 | Ouqvx4);
assign Vcnvx4 = (~(Vuqvx4 & Cvqvx4));
assign Cvqvx4 = (~(Jvqvx4 & hrdata_i[0]));
assign Vuqvx4 = (Qvqvx4 & Xvqvx4);
assign Xvqvx4 = (Ewqvx4 | Abovx4);
assign Qvqvx4 = (~(Hnevx4 & Lwqvx4));
assign Ocnvx4 = (~(Swqvx4 & Zwqvx4));
assign Zwqvx4 = (Gxqvx4 | Nxqvx4);
assign Swqvx4 = (Uxqvx4 & Byqvx4);
assign Byqvx4 = (~(Ouqvx4 & Iyqvx4));
assign Uxqvx4 = (~(Pyqvx4 & F9pvx4));
assign Hcnvx4 = (~(Wyqvx4 & Dzqvx4));
assign Dzqvx4 = (Kzqvx4 | Abovx4);
assign Wyqvx4 = (Rzqvx4 & Yzqvx4);
assign Yzqvx4 = (~(Roevx4 & Lwqvx4));
assign Rzqvx4 = (~(Jvqvx4 & hrdata_i[1]));
assign Acnvx4 = (~(F0rvx4 & M0rvx4));
assign M0rvx4 = (T0rvx4 | Nxqvx4);
assign F0rvx4 = (A1rvx4 & H1rvx4);
assign H1rvx4 = (~(O1rvx4 & Roevx4));
assign A1rvx4 = (~(Pyqvx4 & V1rvx4));
assign V1rvx4 = (!C2rvx4);
assign Tbnvx4 = (~(J2rvx4 & Q2rvx4));
assign Q2rvx4 = (~(X2rvx4 & E3rvx4));
assign J2rvx4 = (L3rvx4 & S3rvx4);
assign S3rvx4 = (~(Bqevx4 & Lwqvx4));
assign L3rvx4 = (~(hrdata_i[2] & Jvqvx4));
assign Mbnvx4 = (~(Z3rvx4 & G4rvx4));
assign G4rvx4 = (~(N4rvx4 & E3rvx4));
assign Z3rvx4 = (U4rvx4 & B5rvx4);
assign B5rvx4 = (~(Lrevx4 & Lwqvx4));
assign U4rvx4 = (~(hrdata_i[3] & Jvqvx4));
assign Fbnvx4 = (~(I5rvx4 & P5rvx4));
assign P5rvx4 = (~(W5rvx4 & E3rvx4));
assign I5rvx4 = (D6rvx4 & K6rvx4);
assign K6rvx4 = (~(Vsevx4 & Lwqvx4));
assign D6rvx4 = (~(Jvqvx4 & hrdata_i[4]));
assign Yanvx4 = (~(R6rvx4 & Y6rvx4));
assign Y6rvx4 = (~(Fuevx4 & Lwqvx4));
assign Lwqvx4 = (~(F7rvx4 & M7rvx4));
assign M7rvx4 = (E3rvx4 | T7rvx4);
assign R6rvx4 = (~(Jvqvx4 & hrdata_i[5]));
assign Ranvx4 = (~(A8rvx4 & H8rvx4));
assign H8rvx4 = (~(Edovx4 & Pvevx4));
assign A8rvx4 = (O8rvx4 & V8rvx4);
assign V8rvx4 = (~(Enh2z4[1] & C9rvx4));
assign O8rvx4 = (~(hrdata_i[6] & Jvqvx4));
assign Kanvx4 = (~(J9rvx4 & Q9rvx4));
assign Q9rvx4 = (~(Edovx4 & Zwevx4));
assign J9rvx4 = (X9rvx4 & Earvx4);
assign Earvx4 = (~(Enh2z4[2] & C9rvx4));
assign X9rvx4 = (~(Jvqvx4 & hrdata_i[7]));
assign Danvx4 = (~(Larvx4 & Sarvx4));
assign Sarvx4 = (~(Edovx4 & Jyevx4));
assign Larvx4 = (Zarvx4 & Gbrvx4);
assign Gbrvx4 = (~(Enh2z4[3] & C9rvx4));
assign Zarvx4 = (~(Jvqvx4 & hrdata_i[8]));
assign W9nvx4 = (~(Nbrvx4 & Ubrvx4));
assign Ubrvx4 = (~(Edovx4 & Tzevx4));
assign Nbrvx4 = (Bcrvx4 & Icrvx4);
assign Icrvx4 = (~(Enh2z4[4] & C9rvx4));
assign Bcrvx4 = (~(Jvqvx4 & hrdata_i[9]));
assign P9nvx4 = (~(Pcrvx4 & Wcrvx4));
assign Wcrvx4 = (~(Edovx4 & D1fvx4));
assign Pcrvx4 = (Ddrvx4 & Kdrvx4);
assign Kdrvx4 = (~(Enh2z4[5] & C9rvx4));
assign Ddrvx4 = (~(hrdata_i[10] & Jvqvx4));
assign I9nvx4 = (~(Rdrvx4 & Ydrvx4));
assign Ydrvx4 = (~(Edovx4 & O2fvx4));
assign Rdrvx4 = (Fervx4 & Mervx4);
assign Mervx4 = (~(Enh2z4[6] & C9rvx4));
assign Fervx4 = (~(hrdata_i[11] & Jvqvx4));
assign B9nvx4 = (~(Tervx4 & Afrvx4));
assign Afrvx4 = (~(Edovx4 & Z3fvx4));
assign Tervx4 = (Hfrvx4 & Ofrvx4);
assign Ofrvx4 = (~(Enh2z4[7] & C9rvx4));
assign Hfrvx4 = (~(Jvqvx4 & hrdata_i[12]));
assign U8nvx4 = (~(Vfrvx4 & Cgrvx4));
assign Cgrvx4 = (~(Edovx4 & K5fvx4));
assign Vfrvx4 = (Jgrvx4 & Qgrvx4);
assign Qgrvx4 = (~(Enh2z4[8] & C9rvx4));
assign C9rvx4 = (Xgrvx4 & Qcovx4);
assign Xgrvx4 = (~(E3rvx4 & Ehrvx4));
assign Ehrvx4 = (~(Lhrvx4 & Shrvx4));
assign Shrvx4 = (Zhrvx4 & Girvx4);
assign Girvx4 = (~(Nirvx4 | Fuevx4));
assign Nirvx4 = (Uirvx4 & Bjrvx4);
assign Bjrvx4 = (~(Ijrvx4 & Roevx4));
assign Ijrvx4 = (Xlevx4 & Pjrvx4);
assign Uirvx4 = (~(Kzqvx4 & Pjrvx4));
assign Pjrvx4 = (Ewqvx4 | Iyqvx4);
assign Iyqvx4 = (!Tnpvx4);
assign Zhrvx4 = (Wjrvx4 & Dkrvx4);
assign Dkrvx4 = (~(Kzqvx4 & Roevx4));
assign Wjrvx4 = (Tnpvx4 | Kkrvx4);
assign Tnpvx4 = (~(Hnevx4 & Xlevx4));
assign Lhrvx4 = (Rkrvx4 & Ykrvx4);
assign Ykrvx4 = (~(N4rvx4 ^ Lrevx4));
assign Rkrvx4 = (Flrvx4 & Mlrvx4);
assign Mlrvx4 = (~(X2rvx4 ^ Bqevx4));
assign Flrvx4 = (Tlrvx4 ^ W5rvx4);
assign Tlrvx4 = (~(Vsevx4 & Xlevx4));
assign Jgrvx4 = (~(Jvqvx4 & hrdata_i[13]));
assign N8nvx4 = (~(Amrvx4 & Hmrvx4));
assign Hmrvx4 = (~(hrdata_i[14] & Jvqvx4));
assign Jvqvx4 = (Omrvx4 & Ueovx4);
assign Omrvx4 = (~(Qcovx4 | Edovx4));
assign Amrvx4 = (~(V6fvx4 & Edovx4));
assign G8nvx4 = (Vmrvx4 | Qcovx4);
assign Vmrvx4 = (F7rvx4 ? Cnrvx4 : G8fvx4);
assign Cnrvx4 = (Ueovx4 & hrdata_i[15]);
assign Z7nvx4 = (!Jnrvx4);
assign Jnrvx4 = (F7rvx4 ? Qcovx4 : Qnrvx4);
assign F7rvx4 = (!Edovx4);
assign Edovx4 = (T7rvx4 & Xnrvx4);
assign Xnrvx4 = (~(Eorvx4 & Lorvx4));
assign Lorvx4 = (~(Wnnvx4 | Cn8vx4));
assign Eorvx4 = (~(Sorvx4 | Zorvx4));
assign Qcovx4 = (!T7rvx4);
assign T7rvx4 = (~(E3rvx4 | Xlevx4));
assign E3rvx4 = (!Abovx4);
assign Qnrvx4 = (~(Gprvx4 & V8evx4));
assign Gprvx4 = (~(Zorvx4 | Wfovx4));
assign S7nvx4 = (~(Nprvx4 & Uprvx4));
assign Uprvx4 = (Bqrvx4 & Iqrvx4);
assign Iqrvx4 = (~(hrdata_i[1] & Vapvx4));
assign Bqrvx4 = (Pqrvx4 & Wqrvx4);
assign Wqrvx4 = (~(Mcfvx4 & Pfovx4));
assign Pqrvx4 = (~(hrdata_i[17] & Qbpvx4));
assign Nprvx4 = (Drrvx4 & Krrvx4);
assign Krrvx4 = (~(Roevx4 & Wfovx4));
assign Drrvx4 = (~(B19vx4 & Geovx4));
assign L7nvx4 = (~(Rrrvx4 & Yrrvx4));
assign Yrrvx4 = (Fsrvx4 & Msrvx4);
assign Msrvx4 = (~(hrdata_i[2] & Vapvx4));
assign Fsrvx4 = (Tsrvx4 & Atrvx4);
assign Atrvx4 = (~(Wdfvx4 & Pfovx4));
assign Tsrvx4 = (~(hrdata_i[18] & Qbpvx4));
assign Rrrvx4 = (Htrvx4 & Otrvx4);
assign Otrvx4 = (~(Bqevx4 & Wfovx4));
assign Htrvx4 = (Vtrvx4 | Scpvx4);
assign E7nvx4 = (~(Curvx4 & Jurvx4));
assign Jurvx4 = (Qurvx4 & Xurvx4);
assign Xurvx4 = (~(hrdata_i[3] & Vapvx4));
assign Qurvx4 = (Evrvx4 & Lvrvx4);
assign Lvrvx4 = (~(Gffvx4 & Pfovx4));
assign Evrvx4 = (~(hrdata_i[19] & Qbpvx4));
assign Curvx4 = (Svrvx4 & Zvrvx4);
assign Zvrvx4 = (~(Lrevx4 & Wfovx4));
assign Svrvx4 = (Gwrvx4 | Scpvx4);
assign X6nvx4 = (~(Nwrvx4 & Uwrvx4));
assign Uwrvx4 = (Bxrvx4 & Ixrvx4);
assign Ixrvx4 = (~(hrdata_i[4] & Vapvx4));
assign Bxrvx4 = (Pxrvx4 & Wxrvx4);
assign Wxrvx4 = (~(Qgfvx4 & Pfovx4));
assign Pxrvx4 = (~(hrdata_i[20] & Qbpvx4));
assign Nwrvx4 = (Dyrvx4 & Kyrvx4);
assign Kyrvx4 = (~(Vsevx4 & Wfovx4));
assign Dyrvx4 = (Ryrvx4 | Scpvx4);
assign Q6nvx4 = (~(Yyrvx4 & Fzrvx4));
assign Fzrvx4 = (Mzrvx4 & Tzrvx4);
assign Tzrvx4 = (~(hrdata_i[5] & Vapvx4));
assign Mzrvx4 = (A0svx4 & H0svx4);
assign H0svx4 = (~(Aifvx4 & Pfovx4));
assign A0svx4 = (~(hrdata_i[21] & Qbpvx4));
assign Yyrvx4 = (O0svx4 & V0svx4);
assign V0svx4 = (~(Fuevx4 & Wfovx4));
assign O0svx4 = (C1svx4 | Scpvx4);
assign J6nvx4 = (~(J1svx4 & Q1svx4));
assign Q1svx4 = (X1svx4 & E2svx4);
assign E2svx4 = (~(hrdata_i[6] & Vapvx4));
assign X1svx4 = (L2svx4 & S2svx4);
assign S2svx4 = (~(Kjfvx4 & Pfovx4));
assign L2svx4 = (~(hrdata_i[22] & Qbpvx4));
assign J1svx4 = (Z2svx4 & G3svx4);
assign G3svx4 = (~(Wfovx4 & Pvevx4));
assign Z2svx4 = (N3svx4 | Scpvx4);
assign C6nvx4 = (~(U3svx4 & B4svx4));
assign B4svx4 = (I4svx4 & P4svx4);
assign P4svx4 = (~(Vapvx4 & hrdata_i[7]));
assign I4svx4 = (W4svx4 & D5svx4);
assign D5svx4 = (~(Ukfvx4 & Pfovx4));
assign W4svx4 = (~(Qbpvx4 & hrdata_i[23]));
assign U3svx4 = (K5svx4 & R5svx4);
assign R5svx4 = (~(Wfovx4 & Zwevx4));
assign K5svx4 = (Y5svx4 | Scpvx4);
assign V5nvx4 = (~(F6svx4 & M6svx4));
assign M6svx4 = (T6svx4 & A7svx4);
assign A7svx4 = (~(Vapvx4 & hrdata_i[8]));
assign T6svx4 = (H7svx4 & O7svx4);
assign O7svx4 = (~(Emfvx4 & Pfovx4));
assign H7svx4 = (~(Qbpvx4 & hrdata_i[24]));
assign F6svx4 = (V7svx4 & C8svx4);
assign C8svx4 = (~(Wfovx4 & Jyevx4));
assign V7svx4 = (J8svx4 | Scpvx4);
assign O5nvx4 = (~(Q8svx4 & X8svx4));
assign X8svx4 = (E9svx4 & L9svx4);
assign L9svx4 = (~(hrdata_i[9] & Vapvx4));
assign E9svx4 = (S9svx4 & Z9svx4);
assign Z9svx4 = (~(Onfvx4 & Pfovx4));
assign S9svx4 = (~(hrdata_i[25] & Qbpvx4));
assign Q8svx4 = (Gasvx4 & Nasvx4);
assign Nasvx4 = (~(Wfovx4 & Tzevx4));
assign Gasvx4 = (Uasvx4 | Scpvx4);
assign H5nvx4 = (~(Bbsvx4 & Ibsvx4));
assign Ibsvx4 = (Pbsvx4 & Wbsvx4);
assign Wbsvx4 = (~(hrdata_i[10] & Vapvx4));
assign Pbsvx4 = (Dcsvx4 & Kcsvx4);
assign Kcsvx4 = (~(Yofvx4 & Pfovx4));
assign Dcsvx4 = (~(hrdata_i[26] & Qbpvx4));
assign Bbsvx4 = (Rcsvx4 & Ycsvx4);
assign Ycsvx4 = (~(Wfovx4 & D1fvx4));
assign Rcsvx4 = (Fdsvx4 | Scpvx4);
assign A5nvx4 = (~(Mdsvx4 & Tdsvx4));
assign Tdsvx4 = (Aesvx4 & Hesvx4);
assign Hesvx4 = (~(hrdata_i[11] & Vapvx4));
assign Aesvx4 = (Oesvx4 & Vesvx4);
assign Vesvx4 = (~(Jqfvx4 & Pfovx4));
assign Oesvx4 = (~(hrdata_i[27] & Qbpvx4));
assign Mdsvx4 = (Cfsvx4 & Jfsvx4);
assign Jfsvx4 = (~(Wfovx4 & O2fvx4));
assign Cfsvx4 = (Qfsvx4 | Scpvx4);
assign T4nvx4 = (~(Xfsvx4 & Egsvx4));
assign Egsvx4 = (Lgsvx4 & Sgsvx4);
assign Sgsvx4 = (~(hrdata_i[12] & Vapvx4));
assign Lgsvx4 = (Zgsvx4 & Ghsvx4);
assign Ghsvx4 = (~(Urfvx4 & Pfovx4));
assign Zgsvx4 = (~(hrdata_i[28] & Qbpvx4));
assign Xfsvx4 = (Nhsvx4 & Uhsvx4);
assign Uhsvx4 = (~(Wfovx4 & Z3fvx4));
assign Nhsvx4 = (Bisvx4 | Scpvx4);
assign M4nvx4 = (~(Iisvx4 & Pisvx4));
assign Pisvx4 = (Wisvx4 & Djsvx4);
assign Djsvx4 = (~(hrdata_i[14] & Vapvx4));
assign Vapvx4 = (Kjsvx4 & Rjsvx4);
assign Rjsvx4 = (~(Neovx4 | Yjsvx4));
assign Kjsvx4 = (~(Xcovx4 | Geovx4));
assign Geovx4 = (!Scpvx4);
assign Wisvx4 = (Fksvx4 & Mksvx4);
assign Mksvx4 = (~(Qufvx4 & Pfovx4));
assign Pfovx4 = (Tksvx4 & Scpvx4);
assign Tksvx4 = (Alsvx4 & Neovx4);
assign Alsvx4 = (~(Hlsvx4 & Olsvx4));
assign Olsvx4 = (Vlsvx4 | V8evx4);
assign Fksvx4 = (~(hrdata_i[30] & Qbpvx4));
assign Qbpvx4 = (Cmsvx4 & Ueovx4);
assign Cmsvx4 = (Yjsvx4 & Scpvx4);
assign Yjsvx4 = (~(Vlsvx4 | Cn8vx4));
assign Iisvx4 = (Jmsvx4 & Qmsvx4);
assign Qmsvx4 = (~(V6fvx4 & Wfovx4));
assign Wfovx4 = (V8evx4 & Scpvx4);
assign Jmsvx4 = (Xmsvx4 | Scpvx4);
assign Scpvx4 = (Ensvx4 & Lnsvx4);
assign Lnsvx4 = (Snsvx4 & Znsvx4);
assign Znsvx4 = (~(Gosvx4 & Nosvx4));
assign Nosvx4 = (~(Uosvx4 & Bpsvx4));
assign Uosvx4 = (Hlsvx4 & Wnnvx4);
assign Snsvx4 = (Ipsvx4 & Z5pvx4);
assign Ensvx4 = (Ppsvx4 & Wpsvx4);
assign F4nvx4 = (S6ovx4 ? hwrite_o : Dqsvx4);
assign S6ovx4 = (Kqsvx4 & Rqsvx4);
assign Rqsvx4 = (Yqsvx4 & Frsvx4);
assign Frsvx4 = (~(Mrsvx4 | haddr_o[28]));
assign Yqsvx4 = (~(W6qvx4 | Trsvx4));
assign Kqsvx4 = (Assvx4 & U5qvx4);
assign Assvx4 = (Hssvx4 & Ppsvx4);
assign Dqsvx4 = (Ossvx4 & Vssvx4);
assign Ossvx4 = (~(Ctsvx4 | Z7hvx4));
assign Y3nvx4 = (~(Jtsvx4 & Qtsvx4));
assign Qtsvx4 = (~(L0i2z4[15] & Xtsvx4));
assign Xtsvx4 = (~(hwdata_o[15] & Zyovx4));
assign Jtsvx4 = (~(hwdata_o[15] & Gzovx4));
assign R3nvx4 = (~(Eusvx4 & Lusvx4));
assign Lusvx4 = (~(L0i2z4[14] & Susvx4));
assign Susvx4 = (~(Zyovx4 & hwdata_o[14]));
assign Eusvx4 = (~(Gzovx4 & hwdata_o[14]));
assign K3nvx4 = (~(Zusvx4 & Gvsvx4));
assign Gvsvx4 = (~(L0i2z4[13] & Nvsvx4));
assign Nvsvx4 = (~(hwdata_o[13] & Zyovx4));
assign Zusvx4 = (~(hwdata_o[13] & Gzovx4));
assign D3nvx4 = (~(Uvsvx4 & Bwsvx4));
assign Bwsvx4 = (~(L0i2z4[12] & Iwsvx4));
assign Iwsvx4 = (~(hwdata_o[12] & Zyovx4));
assign Uvsvx4 = (~(hwdata_o[12] & Gzovx4));
assign W2nvx4 = (~(Pwsvx4 & Wwsvx4));
assign Wwsvx4 = (~(L0i2z4[11] & Dxsvx4));
assign Dxsvx4 = (~(hwdata_o[11] & Zyovx4));
assign Pwsvx4 = (~(hwdata_o[11] & Gzovx4));
assign P2nvx4 = (~(Kxsvx4 & Rxsvx4));
assign Rxsvx4 = (~(L0i2z4[10] & Yxsvx4));
assign Yxsvx4 = (~(hwdata_o[10] & Zyovx4));
assign Kxsvx4 = (~(hwdata_o[10] & Gzovx4));
assign I2nvx4 = (~(Fysvx4 & Mysvx4));
assign Mysvx4 = (~(L0i2z4[9] & Tysvx4));
assign Tysvx4 = (~(hwdata_o[9] & Zyovx4));
assign Fysvx4 = (~(hwdata_o[9] & Gzovx4));
assign B2nvx4 = (~(Azsvx4 & Hzsvx4));
assign Hzsvx4 = (~(L0i2z4[8] & Ozsvx4));
assign Ozsvx4 = (~(hwdata_o[8] & Zyovx4));
assign Azsvx4 = (~(hwdata_o[8] & Gzovx4));
assign U1nvx4 = (~(Vzsvx4 & C0tvx4));
assign C0tvx4 = (~(L0i2z4[7] & J0tvx4));
assign J0tvx4 = (~(hwdata_o[7] & Zyovx4));
assign Vzsvx4 = (~(hwdata_o[7] & Gzovx4));
assign N1nvx4 = (~(Q0tvx4 & X0tvx4));
assign X0tvx4 = (~(L0i2z4[6] & E1tvx4));
assign E1tvx4 = (~(hwdata_o[6] & Zyovx4));
assign Q0tvx4 = (~(hwdata_o[6] & Gzovx4));
assign G1nvx4 = (~(L1tvx4 & S1tvx4));
assign S1tvx4 = (~(L0i2z4[5] & Z1tvx4));
assign Z1tvx4 = (~(hwdata_o[5] & Zyovx4));
assign L1tvx4 = (~(hwdata_o[5] & Gzovx4));
assign Z0nvx4 = (~(G2tvx4 & N2tvx4));
assign N2tvx4 = (~(L0i2z4[4] & U2tvx4));
assign U2tvx4 = (~(hwdata_o[4] & Zyovx4));
assign G2tvx4 = (~(hwdata_o[4] & Gzovx4));
assign S0nvx4 = (~(B3tvx4 & I3tvx4));
assign I3tvx4 = (~(L0i2z4[3] & P3tvx4));
assign P3tvx4 = (~(hwdata_o[3] & Zyovx4));
assign B3tvx4 = (~(hwdata_o[3] & Gzovx4));
assign L0nvx4 = (~(W3tvx4 & D4tvx4));
assign D4tvx4 = (~(L0i2z4[2] & K4tvx4));
assign K4tvx4 = (~(hwdata_o[2] & Zyovx4));
assign W3tvx4 = (~(hwdata_o[2] & Gzovx4));
assign E0nvx4 = (~(R4tvx4 & Y4tvx4));
assign Y4tvx4 = (~(L0i2z4[1] & F5tvx4));
assign F5tvx4 = (~(hwdata_o[1] & Zyovx4));
assign R4tvx4 = (~(hwdata_o[1] & Gzovx4));
assign Gzovx4 = (Zyovx4 & Rgovx4);
assign Zyovx4 = (M5tvx4 & Mf8vx4);
assign Xzmvx4 = (T5tvx4 ? hwdata_o[0] : F2hvx4);
assign Qzmvx4 = (T5tvx4 ? hwdata_o[1] : S0hvx4);
assign T5tvx4 = (A6tvx4 & Mf8vx4);
assign Jzmvx4 = (C5ovx4 ? hwdata_o[0] : Czh2z4[0]);
assign Czmvx4 = (C5ovx4 ? hwdata_o[1] : Czh2z4[1]);
assign Vymvx4 = (C5ovx4 ? hwdata_o[2] : Czh2z4[2]);
assign Oymvx4 = (C5ovx4 ? hwdata_o[3] : Czh2z4[3]);
assign Hymvx4 = (C5ovx4 ? hwdata_o[4] : Czh2z4[4]);
assign Aymvx4 = (C5ovx4 ? hwdata_o[5] : Czh2z4[5]);
assign Txmvx4 = (C5ovx4 ? hwdata_o[6] : Czh2z4[6]);
assign Mxmvx4 = (C5ovx4 ? hwdata_o[7] : Czh2z4[7]);
assign Fxmvx4 = (C5ovx4 ? hwdata_o[8] : Czh2z4[8]);
assign Ywmvx4 = (C5ovx4 ? hwdata_o[9] : Czh2z4[9]);
assign Rwmvx4 = (C5ovx4 ? hwdata_o[10] : Czh2z4[10]);
assign Kwmvx4 = (C5ovx4 ? hwdata_o[11] : Czh2z4[11]);
assign Dwmvx4 = (C5ovx4 ? hwdata_o[12] : Czh2z4[12]);
assign Wvmvx4 = (C5ovx4 ? hwdata_o[13] : Czh2z4[13]);
assign Pvmvx4 = (C5ovx4 ? hwdata_o[14] : Czh2z4[14]);
assign Ivmvx4 = (C5ovx4 ? hwdata_o[15] : Czh2z4[15]);
assign Bvmvx4 = (C5ovx4 ? hwdata_o[16] : Czh2z4[16]);
assign Uumvx4 = (C5ovx4 ? hwdata_o[17] : Czh2z4[17]);
assign Numvx4 = (C5ovx4 ? hwdata_o[18] : Czh2z4[18]);
assign Gumvx4 = (C5ovx4 ? hwdata_o[19] : Czh2z4[19]);
assign Ztmvx4 = (C5ovx4 ? hwdata_o[20] : Czh2z4[20]);
assign Stmvx4 = (C5ovx4 ? hwdata_o[21] : Czh2z4[21]);
assign Ltmvx4 = (C5ovx4 ? hwdata_o[22] : Czh2z4[22]);
assign C5ovx4 = (H6tvx4 & Mf8vx4);
assign Etmvx4 = (~(O6tvx4 & V6tvx4));
assign V6tvx4 = (~(C7tvx4 & Irh2z4[0]));
assign O6tvx4 = (J7tvx4 & Q7tvx4);
assign Q7tvx4 = (~(Iwh2z4[0] & X7tvx4));
assign J7tvx4 = (~(E8tvx4 & Czh2z4[0]));
assign Xsmvx4 = (~(L8tvx4 & S8tvx4));
assign S8tvx4 = (~(C7tvx4 & Irh2z4[1]));
assign L8tvx4 = (Z8tvx4 & G9tvx4);
assign G9tvx4 = (~(Iwh2z4[1] & X7tvx4));
assign Z8tvx4 = (~(E8tvx4 & Czh2z4[1]));
assign Qsmvx4 = (~(N9tvx4 & U9tvx4));
assign U9tvx4 = (~(Irh2z4[2] & C7tvx4));
assign N9tvx4 = (Batvx4 & Iatvx4);
assign Iatvx4 = (~(Iwh2z4[2] & X7tvx4));
assign Batvx4 = (~(E8tvx4 & Czh2z4[2]));
assign Jsmvx4 = (~(Patvx4 & Watvx4));
assign Watvx4 = (~(Irh2z4[3] & C7tvx4));
assign Patvx4 = (Dbtvx4 & Kbtvx4);
assign Kbtvx4 = (~(Iwh2z4[3] & X7tvx4));
assign Dbtvx4 = (~(E8tvx4 & Czh2z4[3]));
assign Csmvx4 = (~(Rbtvx4 & Ybtvx4));
assign Ybtvx4 = (~(C7tvx4 & Irh2z4[4]));
assign Rbtvx4 = (Fctvx4 & Mctvx4);
assign Mctvx4 = (~(Iwh2z4[4] & X7tvx4));
assign Fctvx4 = (~(E8tvx4 & Czh2z4[4]));
assign Vrmvx4 = (~(Tctvx4 & Adtvx4));
assign Adtvx4 = (~(C7tvx4 & Irh2z4[5]));
assign Tctvx4 = (Hdtvx4 & Odtvx4);
assign Odtvx4 = (~(Iwh2z4[5] & X7tvx4));
assign Hdtvx4 = (~(E8tvx4 & Czh2z4[5]));
assign Ormvx4 = (~(Vdtvx4 & Cetvx4));
assign Cetvx4 = (~(Irh2z4[6] & C7tvx4));
assign Vdtvx4 = (Jetvx4 & Qetvx4);
assign Qetvx4 = (~(Iwh2z4[6] & X7tvx4));
assign Jetvx4 = (~(E8tvx4 & Czh2z4[6]));
assign Hrmvx4 = (~(Xetvx4 & Eftvx4));
assign Eftvx4 = (~(C7tvx4 & Irh2z4[7]));
assign Xetvx4 = (Lftvx4 & Sftvx4);
assign Sftvx4 = (~(Iwh2z4[7] & X7tvx4));
assign Lftvx4 = (~(E8tvx4 & Czh2z4[7]));
assign Armvx4 = (~(Zftvx4 & Ggtvx4));
assign Ggtvx4 = (~(C7tvx4 & Irh2z4[8]));
assign Zftvx4 = (Ngtvx4 & Ugtvx4);
assign Ugtvx4 = (~(Iwh2z4[8] & X7tvx4));
assign Ngtvx4 = (~(E8tvx4 & Czh2z4[8]));
assign Tqmvx4 = (~(Bhtvx4 & Ihtvx4));
assign Ihtvx4 = (~(C7tvx4 & Irh2z4[9]));
assign Bhtvx4 = (Phtvx4 & Whtvx4);
assign Whtvx4 = (~(Iwh2z4[9] & X7tvx4));
assign Phtvx4 = (~(E8tvx4 & Czh2z4[9]));
assign Mqmvx4 = (~(Ditvx4 & Kitvx4));
assign Kitvx4 = (~(Irh2z4[10] & C7tvx4));
assign Ditvx4 = (Ritvx4 & Yitvx4);
assign Yitvx4 = (~(Iwh2z4[10] & X7tvx4));
assign Ritvx4 = (~(E8tvx4 & Czh2z4[10]));
assign Fqmvx4 = (~(Fjtvx4 & Mjtvx4));
assign Mjtvx4 = (~(Irh2z4[11] & C7tvx4));
assign Fjtvx4 = (Tjtvx4 & Aktvx4);
assign Aktvx4 = (~(Iwh2z4[11] & X7tvx4));
assign Tjtvx4 = (~(E8tvx4 & Czh2z4[11]));
assign Ypmvx4 = (~(Hktvx4 & Oktvx4));
assign Oktvx4 = (~(C7tvx4 & Irh2z4[12]));
assign Hktvx4 = (Vktvx4 & Cltvx4);
assign Cltvx4 = (~(Iwh2z4[12] & X7tvx4));
assign Vktvx4 = (~(E8tvx4 & Czh2z4[12]));
assign Rpmvx4 = (~(Jltvx4 & Qltvx4));
assign Qltvx4 = (~(C7tvx4 & Irh2z4[13]));
assign Jltvx4 = (Xltvx4 & Emtvx4);
assign Emtvx4 = (~(Iwh2z4[13] & X7tvx4));
assign Xltvx4 = (~(E8tvx4 & Czh2z4[13]));
assign Kpmvx4 = (~(Lmtvx4 & Smtvx4));
assign Smtvx4 = (~(Irh2z4[14] & C7tvx4));
assign Lmtvx4 = (Zmtvx4 & Gntvx4);
assign Gntvx4 = (~(Iwh2z4[14] & X7tvx4));
assign Zmtvx4 = (~(E8tvx4 & Czh2z4[14]));
assign Dpmvx4 = (~(Nntvx4 & Untvx4));
assign Untvx4 = (~(C7tvx4 & Irh2z4[15]));
assign Nntvx4 = (Botvx4 & Iotvx4);
assign Iotvx4 = (~(Iwh2z4[15] & X7tvx4));
assign Botvx4 = (~(E8tvx4 & Czh2z4[15]));
assign Womvx4 = (~(Potvx4 & Wotvx4));
assign Wotvx4 = (~(C7tvx4 & Irh2z4[16]));
assign Potvx4 = (Dptvx4 & Kptvx4);
assign Kptvx4 = (~(Iwh2z4[16] & X7tvx4));
assign Dptvx4 = (~(E8tvx4 & Czh2z4[16]));
assign Pomvx4 = (~(Rptvx4 & Yptvx4));
assign Yptvx4 = (~(C7tvx4 & Irh2z4[17]));
assign Rptvx4 = (Fqtvx4 & Mqtvx4);
assign Mqtvx4 = (~(Iwh2z4[17] & X7tvx4));
assign Fqtvx4 = (~(E8tvx4 & Czh2z4[17]));
assign Iomvx4 = (~(Tqtvx4 & Artvx4));
assign Artvx4 = (~(Irh2z4[18] & C7tvx4));
assign Tqtvx4 = (Hrtvx4 & Ortvx4);
assign Ortvx4 = (~(Iwh2z4[18] & X7tvx4));
assign Hrtvx4 = (~(E8tvx4 & Czh2z4[18]));
assign Bomvx4 = (~(Vrtvx4 & Cstvx4));
assign Cstvx4 = (~(Irh2z4[19] & C7tvx4));
assign Vrtvx4 = (Jstvx4 & Qstvx4);
assign Qstvx4 = (~(Iwh2z4[19] & X7tvx4));
assign Jstvx4 = (~(E8tvx4 & Czh2z4[19]));
assign Unmvx4 = (~(Xstvx4 & Ettvx4));
assign Ettvx4 = (~(C7tvx4 & Irh2z4[20]));
assign Xstvx4 = (Lttvx4 & Sttvx4);
assign Sttvx4 = (~(Iwh2z4[20] & X7tvx4));
assign Lttvx4 = (~(E8tvx4 & Czh2z4[20]));
assign Nnmvx4 = (~(Zttvx4 & Gutvx4));
assign Gutvx4 = (~(C7tvx4 & Irh2z4[21]));
assign Zttvx4 = (Nutvx4 & Uutvx4);
assign Uutvx4 = (~(Iwh2z4[21] & X7tvx4));
assign Nutvx4 = (~(E8tvx4 & Czh2z4[21]));
assign Gnmvx4 = (~(Bvtvx4 & Ivtvx4));
assign Ivtvx4 = (~(Irh2z4[22] & C7tvx4));
assign Bvtvx4 = (Pvtvx4 & Wvtvx4);
assign Wvtvx4 = (~(Iwh2z4[22] & X7tvx4));
assign Pvtvx4 = (~(E8tvx4 & Czh2z4[22]));
assign Zmmvx4 = (~(Dwtvx4 & Kwtvx4));
assign Kwtvx4 = (~(C7tvx4 & Irh2z4[23]));
assign Dwtvx4 = (Rwtvx4 & Ywtvx4);
assign Ywtvx4 = (~(Iwh2z4[23] & X7tvx4));
assign X7tvx4 = (Fxtvx4 & Mxtvx4);
assign Fxtvx4 = (~(C7tvx4 | Txtvx4));
assign Rwtvx4 = (~(E8tvx4 & Czh2z4[23]));
assign E8tvx4 = (~(Aytvx4 | Mxtvx4));
assign Mxtvx4 = (Hytvx4 | Irh2z4[0]);
assign Hytvx4 = (!Oytvx4);
assign Aytvx4 = (C7tvx4 | Txtvx4);
assign C7tvx4 = (~(F2hvx4 | Txtvx4));
assign Smmvx4 = (Vytvx4 ? hwdata_o[6] : Zuh2z4[24]);
assign Lmmvx4 = (Vytvx4 ? hwdata_o[7] : Zuh2z4[25]);
assign Emmvx4 = (Vytvx4 ? hwdata_o[14] : Zuh2z4[26]);
assign Xlmvx4 = (Vytvx4 ? hwdata_o[15] : Zuh2z4[27]);
assign Qlmvx4 = (Vytvx4 ? hwdata_o[22] : Zuh2z4[28]);
assign Jlmvx4 = (Vytvx4 ? V4ovx4 : Zuh2z4[29]);
assign Clmvx4 = (Vytvx4 ? hwdata_o[30] : Zuh2z4[30]);
assign Vkmvx4 = (Vytvx4 ? Cztvx4 : Zuh2z4[31]);
assign Vytvx4 = (Jztvx4 & Mf8vx4);
assign Okmvx4 = (Qztvx4 ? hwdata_o[6] : Zuh2z4[16]);
assign Hkmvx4 = (Qztvx4 ? hwdata_o[7] : Zuh2z4[17]);
assign Akmvx4 = (Qztvx4 ? hwdata_o[14] : Zuh2z4[18]);
assign Tjmvx4 = (Qztvx4 ? hwdata_o[15] : Zuh2z4[19]);
assign Mjmvx4 = (Qztvx4 ? hwdata_o[22] : Zuh2z4[20]);
assign Fjmvx4 = (Qztvx4 ? V4ovx4 : Zuh2z4[21]);
assign Yimvx4 = (Qztvx4 ? hwdata_o[30] : Zuh2z4[22]);
assign Rimvx4 = (Qztvx4 ? Cztvx4 : Zuh2z4[23]);
assign Qztvx4 = (Xztvx4 & Mf8vx4);
assign Xztvx4 = (!E0uvx4);
assign Kimvx4 = (L0uvx4 ? hwdata_o[6] : Zuh2z4[8]);
assign Dimvx4 = (L0uvx4 ? hwdata_o[7] : Zuh2z4[9]);
assign Whmvx4 = (L0uvx4 ? hwdata_o[14] : Zuh2z4[10]);
assign Phmvx4 = (L0uvx4 ? hwdata_o[15] : Zuh2z4[11]);
assign Ihmvx4 = (L0uvx4 ? hwdata_o[22] : Zuh2z4[12]);
assign Bhmvx4 = (L0uvx4 ? V4ovx4 : Zuh2z4[13]);
assign Ugmvx4 = (L0uvx4 ? hwdata_o[30] : Zuh2z4[14]);
assign Ngmvx4 = (L0uvx4 ? Cztvx4 : Zuh2z4[15]);
assign L0uvx4 = (S0uvx4 & Mf8vx4);
assign Ggmvx4 = (Z0uvx4 ? hwdata_o[6] : Zuh2z4[0]);
assign Zfmvx4 = (Z0uvx4 ? hwdata_o[7] : Zuh2z4[1]);
assign Sfmvx4 = (Z0uvx4 ? hwdata_o[14] : Zuh2z4[2]);
assign Lfmvx4 = (Z0uvx4 ? hwdata_o[15] : Zuh2z4[3]);
assign Efmvx4 = (Z0uvx4 ? hwdata_o[22] : Zuh2z4[4]);
assign Xemvx4 = (Z0uvx4 ? V4ovx4 : Zuh2z4[5]);
assign Qemvx4 = (Z0uvx4 ? hwdata_o[30] : Zuh2z4[6]);
assign Jemvx4 = (Z0uvx4 ? Cztvx4 : Zuh2z4[7]);
assign Z0uvx4 = (G1uvx4 & Mf8vx4);
assign G1uvx4 = (!N1uvx4);
assign Cemvx4 = (U1uvx4 ? hwdata_o[4] : Vogvx4);
assign Vdmvx4 = (U1uvx4 ? hwdata_o[2] : Nngvx4);
assign Odmvx4 = (U1uvx4 ? hwdata_o[1] : Eg8vx4);
assign U1uvx4 = (B2uvx4 & Mf8vx4);
assign Hdmvx4 = (I2uvx4 ? Uth2z4[0] : hwdata_o[30]);
assign Admvx4 = (I2uvx4 ? Uth2z4[1] : Cztvx4);
assign I2uvx4 = (~(P2uvx4 & Mf8vx4));
assign Tcmvx4 = (W2uvx4 ? hwdata_o[22] : Psh2z4[0]);
assign Mcmvx4 = (W2uvx4 ? V4ovx4 : Psh2z4[1]);
assign Fcmvx4 = (W2uvx4 ? hwdata_o[30] : Txh2z4[0]);
assign Ybmvx4 = (W2uvx4 ? Cztvx4 : Txh2z4[1]);
assign W2uvx4 = (D3uvx4 & Mf8vx4);
assign D3uvx4 = (!K3uvx4);
assign Rbmvx4 = (~(R3uvx4 & Y3uvx4));
assign Y3uvx4 = (~(F4uvx4 & Izgvx4));
assign F4uvx4 = (~(M4uvx4 | Txtvx4));
assign Txtvx4 = (~(T4uvx4 | Ctsvx4));
assign M4uvx4 = (~(A5uvx4 | Mf8vx4));
assign R3uvx4 = (~(H5uvx4 & Oytvx4));
assign Kbmvx4 = (O5uvx4 & irq_i[15]);
assign O5uvx4 = (V5uvx4 & C6uvx4);
assign C6uvx4 = (~(J6uvx4 & Q6uvx4));
assign V5uvx4 = (~(X6uvx4 & E7uvx4));
assign E7uvx4 = (hwdata_o[15] | L7uvx4);
assign X6uvx4 = (S7uvx4 & Y9ovx4);
assign S7uvx4 = (~(Z7uvx4 & G8uvx4));
assign Dbmvx4 = (N8uvx4 & irq_i[13]);
assign N8uvx4 = (U8uvx4 & B9uvx4);
assign B9uvx4 = (~(I9uvx4 & P9uvx4));
assign U8uvx4 = (~(W9uvx4 & Dauvx4));
assign Dauvx4 = (hwdata_o[13] | L7uvx4);
assign W9uvx4 = (Kauvx4 & Y9ovx4);
assign Kauvx4 = (~(Rauvx4 & Yauvx4));
assign Wamvx4 = (~(Fbuvx4 & Mbuvx4));
assign Mbuvx4 = (~(vis_ipsr_o[5] & Tbuvx4));
assign Fbuvx4 = (Acuvx4 & Hcuvx4);
assign Hcuvx4 = (~(Fuevx4 & O1rvx4));
assign Acuvx4 = (~(Pyqvx4 & Ocuvx4));
assign Ocuvx4 = (!Vcuvx4);
assign Pamvx4 = (~(Cduvx4 & Jduvx4));
assign Jduvx4 = (~(vis_ipsr_o[4] & Tbuvx4));
assign Tbuvx4 = (!Nxqvx4);
assign Cduvx4 = (Qduvx4 & Xduvx4);
assign Xduvx4 = (~(Vsevx4 & O1rvx4));
assign Qduvx4 = (~(Pyqvx4 & Eeuvx4));
assign Eeuvx4 = (!Leuvx4);
assign Iamvx4 = (Seuvx4 & irq_i[3]);
assign Seuvx4 = (Zeuvx4 & Gfuvx4);
assign Gfuvx4 = (~(Nfuvx4 & Ufuvx4));
assign Zeuvx4 = (~(Bguvx4 & Iguvx4));
assign Iguvx4 = (D9ovx4 | Pguvx4);
assign Bguvx4 = (Wguvx4 & Y9ovx4);
assign Wguvx4 = (Dhuvx4 | hwdata_o[3]);
assign Dhuvx4 = (~(Maovx4 | Khuvx4));
assign Bamvx4 = (Rhuvx4 & irq_i[2]);
assign Rhuvx4 = (Yhuvx4 & Fiuvx4);
assign Fiuvx4 = (~(Miuvx4 & Tiuvx4));
assign Yhuvx4 = (~(Ajuvx4 & Hjuvx4));
assign Hjuvx4 = (hwdata_o[2] | L7uvx4);
assign Ajuvx4 = (Ojuvx4 & Y9ovx4);
assign Ojuvx4 = (~(Vjuvx4 & Ckuvx4));
assign U9mvx4 = (~(Jkuvx4 & Qkuvx4));
assign Qkuvx4 = (Xkuvx4 | Nxqvx4);
assign Jkuvx4 = (Eluvx4 & Lluvx4);
assign Lluvx4 = (~(Bqevx4 & O1rvx4));
assign Eluvx4 = (~(Pyqvx4 & Sluvx4));
assign Sluvx4 = (!Zluvx4);
assign N9mvx4 = (Gmuvx4 & irq_i[7]);
assign Gmuvx4 = (Nmuvx4 & Umuvx4);
assign Umuvx4 = (~(Bnuvx4 & Inuvx4));
assign Nmuvx4 = (~(Pnuvx4 & Wnuvx4));
assign Wnuvx4 = (Douvx4 | D9ovx4);
assign Pnuvx4 = (Kouvx4 & Y9ovx4);
assign Kouvx4 = (~(Rouvx4 & Youvx4));
assign Rouvx4 = (Maovx4 | Fpuvx4);
assign G9mvx4 = (Mpuvx4 & irq_i[6]);
assign Mpuvx4 = (Tpuvx4 & Aquvx4);
assign Aquvx4 = (~(Hquvx4 & Oquvx4));
assign Tpuvx4 = (~(Vquvx4 & Cruvx4));
assign Cruvx4 = (D9ovx4 | Jruvx4);
assign Vquvx4 = (Qruvx4 & Y9ovx4);
assign Qruvx4 = (Xruvx4 | hwdata_o[6]);
assign Xruvx4 = (~(Maovx4 | Esuvx4));
assign Z8mvx4 = (Lsuvx4 & irq_i[5]);
assign Lsuvx4 = (Ssuvx4 & Zsuvx4);
assign Zsuvx4 = (~(Gtuvx4 & Ntuvx4));
assign Ssuvx4 = (~(Utuvx4 & Buuvx4));
assign Buuvx4 = (D9ovx4 | Iuuvx4);
assign Utuvx4 = (Puuvx4 & Y9ovx4);
assign Puuvx4 = (~(Wuuvx4 & Dvuvx4));
assign Wuuvx4 = (Maovx4 | Kvuvx4);
assign S8mvx4 = (Rvuvx4 & irq_i[4]);
assign Rvuvx4 = (Yvuvx4 & Fwuvx4);
assign Fwuvx4 = (~(Mwuvx4 & Twuvx4));
assign Yvuvx4 = (~(Axuvx4 & Hxuvx4));
assign Hxuvx4 = (D9ovx4 | Oxuvx4);
assign Axuvx4 = (Vxuvx4 & Y9ovx4);
assign Vxuvx4 = (~(Cyuvx4 & Jyuvx4));
assign Cyuvx4 = (Maovx4 | Qyuvx4);
assign L8mvx4 = (~(Xyuvx4 & Ezuvx4));
assign Ezuvx4 = (Lzuvx4 | Nxqvx4);
assign Xyuvx4 = (Szuvx4 & Zzuvx4);
assign Zzuvx4 = (~(Lrevx4 & O1rvx4));
assign O1rvx4 = (Ouqvx4 & Xlevx4);
assign Ouqvx4 = (Nxqvx4 & G0vvx4);
assign G0vvx4 = (Huqvx4 | Auqvx4);
assign Szuvx4 = (~(Pyqvx4 & N0vvx4));
assign N0vvx4 = (!U0vvx4);
assign Pyqvx4 = (Nxqvx4 & B1vvx4);
assign E8mvx4 = (I1vvx4 & P1vvx4);
assign P1vvx4 = (W1vvx4 & D2vvx4);
assign W1vvx4 = (~(K2vvx4 & R2vvx4));
assign I1vvx4 = (nmi_i & Y2vvx4);
assign Y2vvx4 = (~(L7uvx4 & F3vvx4));
assign X7mvx4 = (~(M3vvx4 & T3vvx4));
assign T3vvx4 = (A4vvx4 | H4vvx4);
assign H4vvx4 = (C5vvx4 ? V4vvx4 : O4vvx4);
assign V4vvx4 = (~(Mtqvx4 & F3vvx4));
assign A4vvx4 = (~(J5vvx4 & Dmgvx4));
assign M3vvx4 = (~(Ul8vx4 & Gosvx4));
assign Q7mvx4 = (~(Q5vvx4 & X5vvx4));
assign X5vvx4 = (~(Krgvx4 & E6vvx4));
assign E6vvx4 = (~(L6vvx4 & vis_ipsr_o[0]));
assign L6vvx4 = (~(Vbovx4 | S6vvx4));
assign J7mvx4 = (Z6vvx4 & irq_i[11]);
assign Z6vvx4 = (G7vvx4 & N7vvx4);
assign N7vvx4 = (~(U7vvx4 & B8vvx4));
assign G7vvx4 = (~(I8vvx4 & P8vvx4));
assign P8vvx4 = (hwdata_o[11] | L7uvx4);
assign I8vvx4 = (W8vvx4 & Y9ovx4);
assign W8vvx4 = (~(D9vvx4 & K9vvx4));
assign C7mvx4 = (R9vvx4 & irq_i[10]);
assign R9vvx4 = (Y9vvx4 & Favvx4);
assign Favvx4 = (~(Mavvx4 & Tavvx4));
assign Y9vvx4 = (~(Abvvx4 & Hbvvx4));
assign Hbvvx4 = (hwdata_o[10] | L7uvx4);
assign Abvvx4 = (Obvvx4 & Y9ovx4);
assign Obvvx4 = (~(Vbvvx4 & Ccvvx4));
assign V6mvx4 = (Jcvvx4 & irq_i[9]);
assign Jcvvx4 = (Qcvvx4 & Xcvvx4);
assign Xcvvx4 = (~(Edvvx4 & Ldvvx4));
assign Qcvvx4 = (~(Sdvvx4 & Zdvvx4));
assign Zdvvx4 = (hwdata_o[9] | L7uvx4);
assign Sdvvx4 = (Gevvx4 & Y9ovx4);
assign Gevvx4 = (~(Nevvx4 & Uevvx4));
assign O6mvx4 = (Bfvvx4 & irq_i[8]);
assign Bfvvx4 = (Ifvvx4 & Pfvvx4);
assign Pfvvx4 = (~(Wfvvx4 & Dgvvx4));
assign Ifvvx4 = (~(Kgvvx4 & Rgvvx4));
assign Rgvvx4 = (hwdata_o[8] | L7uvx4);
assign Kgvvx4 = (Ygvvx4 & Y9ovx4);
assign Ygvvx4 = (~(Fhvvx4 & Mhvvx4));
assign H6mvx4 = (~(Thvvx4 & Aivvx4));
assign Aivvx4 = (~(Wtgvx4 & Hivvx4));
assign Hivvx4 = (Oivvx4 | Vbovx4);
assign Thvvx4 = (Vivvx4 | Cjvvx4);
assign A6mvx4 = (Jjvvx4 & irq_i[12]);
assign Jjvvx4 = (Qjvvx4 & Xjvvx4);
assign Xjvvx4 = (~(Ekvvx4 & Lkvvx4));
assign Qjvvx4 = (~(Skvvx4 & Zkvvx4));
assign Zkvvx4 = (hwdata_o[12] | L7uvx4);
assign Skvvx4 = (Glvvx4 & Y9ovx4);
assign Glvvx4 = (~(Nlvvx4 & Ulvvx4));
assign T5mvx4 = (~(Bmvvx4 & Imvvx4));
assign Imvvx4 = (~(Pmvvx4 & hwdata_o[28]));
assign Bmvvx4 = (~(Wmvvx4 & Qsgvx4));
assign Wmvvx4 = (Dnvvx4 & Knvvx4);
assign Knvvx4 = (~(Pmvvx4 & hwdata_o[27]));
assign Dnvvx4 = (Rnvvx4 | Vbovx4);
assign M5mvx4 = (~(Ynvvx4 & Fovvx4));
assign Fovvx4 = (~(Movvx4 & R3hvx4));
assign Movvx4 = (Tovvx4 & Apvvx4);
assign Apvvx4 = (~(Pmvvx4 & hwdata_o[25]));
assign Tovvx4 = (Hpvvx4 | Vbovx4);
assign F5mvx4 = (~(Opvvx4 & Vpvvx4));
assign Vpvvx4 = (~(Cqvvx4 & Dmgvx4));
assign Cqvvx4 = (Jqvvx4 & C5vvx4);
assign Jqvvx4 = (~(Qqvvx4 & Xqvvx4));
assign Xqvvx4 = (~(Ervvx4 & Lrvvx4));
assign Ervvx4 = (J5vvx4 & Mtqvx4);
assign Qqvvx4 = (~(Srvvx4 & Nxqvx4));
assign Nxqvx4 = (~(Ccovx4 | Mtqvx4));
assign Srvvx4 = (~(Zrvvx4 | vis_pc_o[1]));
assign Opvvx4 = (~(Mk8vx4 & Gosvx4));
assign Gosvx4 = (~(Cn8vx4 & hready_i));
assign Y4mvx4 = (Gsvvx4 & irq_i[1]);
assign Gsvvx4 = (Nsvvx4 & Usvvx4);
assign Usvvx4 = (~(Btvvx4 & Itvvx4));
assign Nsvvx4 = (~(Ptvvx4 & Wtvvx4));
assign Wtvvx4 = (hwdata_o[1] | L7uvx4);
assign Ptvvx4 = (Duvvx4 & Y9ovx4);
assign Duvvx4 = (~(Kuvvx4 & Ruvvx4));
assign R4mvx4 = (Yuvvx4 & irq_i[14]);
assign Yuvvx4 = (Fvvvx4 & Mvvvx4);
assign Mvvvx4 = (~(Tvvvx4 & Awvvx4));
assign Fvvvx4 = (~(Hwvvx4 & Owvvx4));
assign Owvvx4 = (L7uvx4 | hwdata_o[14]);
assign Hwvvx4 = (Vwvvx4 & Y9ovx4);
assign Y9ovx4 = (D9ovx4 | L7uvx4);
assign Vwvvx4 = (~(Cxvvx4 & Jxvvx4));
assign K4mvx4 = (~(Qxvvx4 & Xxvvx4));
assign Xxvvx4 = (Eyvvx4 & Lyvvx4);
assign Lyvvx4 = (R1pvx4 | Fvovx4);
assign Fvovx4 = (Syvvx4 & Zyvvx4);
assign Zyvvx4 = (~(Gzvvx4 & Qrnvx4));
assign Syvvx4 = (Nzvvx4 & Uzvvx4);
assign Uzvvx4 = (~(B0wvx4 & Mrsvx4));
assign B0wvx4 = (I0wvx4 & Bnnvx4);
assign Bnnvx4 = (P0wvx4 | Vlsvx4);
assign P0wvx4 = (Zorvx4 | W0wvx4);
assign I0wvx4 = (~(W0wvx4 & D1wvx4));
assign D1wvx4 = (Vlsvx4 | Zorvx4);
assign W0wvx4 = (~(Wnnvx4 ^ Pnnvx4));
assign Nzvvx4 = (~(Dmh2z4[2] & K1wvx4));
assign Eyvvx4 = (~(P0pvx4 & vis_ipsr_o[2]));
assign Qxvvx4 = (R1wvx4 & Y1wvx4);
assign Y1wvx4 = (~(W0pvx4 & vis_pc_o[1]));
assign R1wvx4 = (~(E1dvx4 & F2pvx4));
assign D4mvx4 = (~(F2wvx4 & M2wvx4));
assign M2wvx4 = (~(Kycvx4 & F2pvx4));
assign F2wvx4 = (T2wvx4 & A3wvx4);
assign A3wvx4 = (~(H3wvx4 & O3wvx4));
assign O3wvx4 = (~(V3wvx4 & C4wvx4));
assign C4wvx4 = (~(vis_tbit_o & J4wvx4));
assign J4wvx4 = (Q4wvx4 | X4wvx4);
assign X4wvx4 = (E5wvx4 & L5wvx4);
assign E5wvx4 = (~(Uasvx4 | J8svx4));
assign T2wvx4 = (~(P0pvx4 & vis_ipsr_o[0]));
assign W3mvx4 = (~(S5wvx4 & Z5wvx4));
assign S5wvx4 = (U6wvx4 ? N6wvx4 : G6wvx4);
assign N6wvx4 = (B7wvx4 & I7wvx4);
assign I7wvx4 = (P7wvx4 | Y5svx4);
assign B7wvx4 = (W7wvx4 & D8wvx4);
assign D8wvx4 = (~(Uz8vx4 & K8wvx4));
assign W7wvx4 = (~(Y99vx4 & R8wvx4));
assign P3mvx4 = (~(Y8wvx4 & F9wvx4));
assign F9wvx4 = (~(U6wvx4 & M9wvx4));
assign M9wvx4 = (~(T9wvx4 & Aawvx4));
assign Aawvx4 = (P7wvx4 | J8svx4);
assign T9wvx4 = (Hawvx4 & Oawvx4);
assign Oawvx4 = (~(B19vx4 & K8wvx4));
assign Hawvx4 = (~(Fb9vx4 & R8wvx4));
assign Y8wvx4 = (Vawvx4 & Z5wvx4);
assign Vawvx4 = (~(Su9vx4 & Cbwvx4));
assign Cbwvx4 = (~(U6wvx4 & Jbwvx4));
assign Jbwvx4 = (~(Ot9vx4 & Qbwvx4));
assign I3mvx4 = (~(Xbwvx4 & Ecwvx4));
assign Ecwvx4 = (Lcwvx4 & Z5wvx4);
assign Lcwvx4 = (~(Wv9vx4 & Scwvx4));
assign Scwvx4 = (~(U6wvx4 & Zcwvx4));
assign Zcwvx4 = (~(Su9vx4 & Qbwvx4));
assign Xbwvx4 = (Gdwvx4 & Ndwvx4);
assign Ndwvx4 = (~(U6wvx4 & Udwvx4));
assign Udwvx4 = (~(Bewvx4 & Iewvx4));
assign Iewvx4 = (P7wvx4 | Uasvx4);
assign Bewvx4 = (Pewvx4 & Wewvx4);
assign Wewvx4 = (~(I29vx4 & K8wvx4));
assign K8wvx4 = (~(Dfwvx4 & Kfwvx4));
assign Kfwvx4 = (Rfwvx4 & Yfwvx4);
assign Yfwvx4 = (~(Fgwvx4 & Mgwvx4));
assign Fgwvx4 = (Tgwvx4 & O4ovx4);
assign Tgwvx4 = (Ahwvx4 | Q4wvx4);
assign Rfwvx4 = (~(Hhwvx4 & Ohwvx4));
assign Hhwvx4 = (~(Bisvx4 | Mc9vx4));
assign Dfwvx4 = (Vhwvx4 & Ciwvx4);
assign Pewvx4 = (~(Mc9vx4 & R8wvx4));
assign R8wvx4 = (~(Jiwvx4 & Qiwvx4));
assign Qiwvx4 = (Xiwvx4 & Ejwvx4);
assign Xiwvx4 = (~(Ljwvx4 & Sjwvx4));
assign Ljwvx4 = (~(Zjwvx4 | Mj8vx4));
assign Jiwvx4 = (Gkwvx4 & Nkwvx4);
assign Nkwvx4 = (~(Ohwvx4 & Ukwvx4));
assign Ukwvx4 = (Bisvx4 | Blwvx4);
assign Gdwvx4 = (~(Ilwvx4 & Qbwvx4));
assign B3mvx4 = (~(Plwvx4 & Wlwvx4));
assign Wlwvx4 = (U6wvx4 ? Kmwvx4 : Dmwvx4);
assign Kmwvx4 = (Rmwvx4 & Ymwvx4);
assign Ymwvx4 = (Fnwvx4 & Mnwvx4);
assign Mnwvx4 = (~(Tnwvx4 & Blwvx4));
assign Fnwvx4 = (Ejwvx4 | Qfsvx4);
assign Ejwvx4 = (~(Aowvx4 & O4ovx4));
assign Aowvx4 = (Howvx4 | Oowvx4);
assign Rmwvx4 = (Vowvx4 & Cpwvx4);
assign Cpwvx4 = (Gwrvx4 | Vhwvx4);
assign Vhwvx4 = (Jpwvx4 & Qpwvx4);
assign Jpwvx4 = (~(Tnwvx4 & Xpwvx4));
assign Xpwvx4 = (Eqwvx4 & Lqwvx4);
assign Eqwvx4 = (Uasvx4 | Qfsvx4);
assign Tnwvx4 = (Ohwvx4 & Cf9vx4);
assign Vowvx4 = (P7wvx4 | Fdsvx4);
assign Plwvx4 = (Sqwvx4 & Z5wvx4);
assign Z5wvx4 = (~(U6wvx4 & Zqwvx4));
assign Zqwvx4 = (~(Grwvx4 & Nrwvx4));
assign Grwvx4 = (Urwvx4 & Bswvx4);
assign Urwvx4 = (~(Iswvx4 & Ukpvx4));
assign Iswvx4 = (Pswvx4 & R89vx4);
assign U6wvx4 = (Wswvx4 & hready_i);
assign Wswvx4 = (~(Dtwvx4 & Ktwvx4));
assign Ktwvx4 = (Rtwvx4 & Ytwvx4);
assign Ytwvx4 = (Fuwvx4 & Muwvx4);
assign Muwvx4 = (Tuwvx4 & Avwvx4);
assign Fuwvx4 = (~(Hvwvx4 | Ovwvx4));
assign Rtwvx4 = (Vvwvx4 & Cwwvx4);
assign Cwwvx4 = (~(B1vvx4 & Jwwvx4));
assign Vvwvx4 = (Qwwvx4 & Xwwvx4);
assign Xwwvx4 = (~(Exwvx4 & Lxwvx4));
assign Exwvx4 = (Sxwvx4 & J8svx4);
assign Sxwvx4 = (~(Lqwvx4 & Zxwvx4));
assign Zxwvx4 = (Gywvx4 | Fdsvx4);
assign Gywvx4 = (!Nywvx4);
assign Qwwvx4 = (~(Uywvx4 & Bzwvx4));
assign Uywvx4 = (~(Izwvx4 | Aj9vx4));
assign Dtwvx4 = (Pzwvx4 & Wzwvx4);
assign Wzwvx4 = (D0xvx4 & K0xvx4);
assign K0xvx4 = (R0xvx4 & Y0xvx4);
assign Y0xvx4 = (F1xvx4 | M1xvx4);
assign R0xvx4 = (~(T1xvx4 & A2xvx4));
assign D0xvx4 = (H2xvx4 & O2xvx4);
assign O2xvx4 = (V2xvx4 | Xmsvx4);
assign V2xvx4 = (!Oowvx4);
assign Pzwvx4 = (C3xvx4 & J3xvx4);
assign C3xvx4 = (Q3xvx4 & X3xvx4);
assign Sqwvx4 = (~(E4xvx4 & Qbwvx4));
assign Qbwvx4 = (~(Zrvvx4 & L4xvx4));
assign L4xvx4 = (~(Ilpvx4 & S4xvx4));
assign U2mvx4 = (Rfpvx4 ? Z4xvx4 : Qm9vx4);
assign Z4xvx4 = (~(G5xvx4 & N5xvx4));
assign N5xvx4 = (U5xvx4 & B6xvx4);
assign B6xvx4 = (I6xvx4 & Hhpvx4);
assign Hhpvx4 = (~(P6xvx4 & W6xvx4));
assign W6xvx4 = (~(D7xvx4 & K7xvx4));
assign D7xvx4 = (Vtrvx4 | Efgvx4);
assign I6xvx4 = (~(R7xvx4 & Xipvx4));
assign R7xvx4 = (Y7xvx4 ^ F8xvx4);
assign U5xvx4 = (M8xvx4 & T8xvx4);
assign T8xvx4 = (~(A9xvx4 & Vopvx4));
assign A9xvx4 = (Qm9vx4 ^ H9xvx4);
assign M8xvx4 = (~(Zpqvx4 & B19vx4));
assign G5xvx4 = (O9xvx4 & V9xvx4);
assign V9xvx4 = (Caxvx4 & Jaxvx4);
assign Jaxvx4 = (~(Bqevx4 & Irqvx4));
assign Caxvx4 = (~(Y99vx4 & Mnpvx4));
assign Mnpvx4 = (~(Qaxvx4 & Xaxvx4));
assign O9xvx4 = (Ebxvx4 & Lbxvx4);
assign Lbxvx4 = (~(I29vx4 & Rmpvx4));
assign Ebxvx4 = (~(Dsqvx4 & R89vx4));
assign N2mvx4 = (Rfpvx4 ? Sbxvx4 : Un9vx4);
assign Rfpvx4 = (Zbxvx4 & hready_i);
assign Zbxvx4 = (~(Gcxvx4 & Ncxvx4));
assign Ncxvx4 = (Ucxvx4 & Bdxvx4);
assign Bdxvx4 = (Idxvx4 & Pdxvx4);
assign Pdxvx4 = (~(Wdxvx4 & Dexvx4));
assign Dexvx4 = (~(O4ovx4 & Kexvx4));
assign Kexvx4 = (Zrvvx4 | Rexvx4);
assign Idxvx4 = (Yexvx4 & Ffxvx4);
assign Yexvx4 = (~(Mfxvx4 & Tfxvx4));
assign Tfxvx4 = (!Agxvx4);
assign Mfxvx4 = (~(Hgxvx4 | U9gvx4));
assign Ucxvx4 = (Ogxvx4 & Vgxvx4);
assign Vgxvx4 = (Chxvx4 | Jhxvx4);
assign Ogxvx4 = (~(Hvwvx4 & Mc9vx4));
assign Hvwvx4 = (Qhxvx4 & Xhxvx4);
assign Qhxvx4 = (~(Ho8vx4 | Sh9vx4));
assign Gcxvx4 = (Eixvx4 & Lixvx4);
assign Lixvx4 = (Sixvx4 & Zixvx4);
assign Zixvx4 = (Agqvx4 | Gjxvx4);
assign Sixvx4 = (Njxvx4 | Ujxvx4);
assign Eixvx4 = (Bkxvx4 & Ikxvx4);
assign Ikxvx4 = (~(Pkxvx4 & Wkxvx4));
assign Sbxvx4 = (~(Dlxvx4 & Klxvx4));
assign Klxvx4 = (Rlxvx4 & Ylxvx4);
assign Ylxvx4 = (Fmxvx4 & Mmxvx4);
assign Mmxvx4 = (~(Tmxvx4 & Vopvx4));
assign Tmxvx4 = (~(Un9vx4 ^ Anxvx4));
assign Fmxvx4 = (Hnxvx4 & Bswvx4);
assign Hnxvx4 = (~(Onxvx4 & Xipvx4));
assign Xipvx4 = (~(Vnxvx4 & Coxvx4));
assign Coxvx4 = (~(Joxvx4 & Qoxvx4));
assign Joxvx4 = (Ukpvx4 & Aj9vx4);
assign Vnxvx4 = (~(Xoxvx4 & Ohwvx4));
assign Xoxvx4 = (~(Epxvx4 | Fdsvx4));
assign Onxvx4 = (~(Lpxvx4 & Spxvx4));
assign Spxvx4 = (~(Y7xvx4 & F8xvx4));
assign F8xvx4 = (Zpxvx4 ^ Gqxvx4);
assign Y7xvx4 = (Coqvx4 & Joqvx4);
assign Joqvx4 = (Nqxvx4 ^ Uqxvx4);
assign Coqvx4 = (Ejpvx4 & Ljpvx4);
assign Ljpvx4 = (~(Brxvx4 ^ Y5svx4));
assign Lpxvx4 = (~(Gqxvx4 & Zpxvx4));
assign Zpxvx4 = (~(Irxvx4 ^ Prxvx4));
assign Prxvx4 = (Wrxvx4 & Dsxvx4);
assign Dsxvx4 = (~(Ksxvx4 & Rsxvx4));
assign Ksxvx4 = (~(N3svx4 | Ysxvx4));
assign Irxvx4 = (~(Ftxvx4 & Mtxvx4));
assign Mtxvx4 = (Ttxvx4 | Auxvx4);
assign Ftxvx4 = (Huxvx4 | Ouxvx4);
assign Gqxvx4 = (Uqxvx4 & Nqxvx4);
assign Nqxvx4 = (~(Vuxvx4 ^ Rsxvx4));
assign Rsxvx4 = (Wrxvx4 & Cvxvx4);
assign Cvxvx4 = (Jvxvx4 | Qvxvx4);
assign Wrxvx4 = (~(Qvxvx4 & Jvxvx4));
assign Jvxvx4 = (Ouxvx4 ^ Huxvx4);
assign Huxvx4 = (~(W49vx4 & Xvxvx4));
assign Ouxvx4 = (~(Ttxvx4 ^ Auxvx4));
assign Auxvx4 = (~(Ewxvx4 | Lwxvx4));
assign Ewxvx4 = (I29vx4 & Swxvx4);
assign Ttxvx4 = (~(P39vx4 & Zwxvx4));
assign Qvxvx4 = (D69vx4 & Gxxvx4);
assign Vuxvx4 = (N3svx4 | Ysxvx4);
assign Uqxvx4 = (R89vx4 & Brxvx4);
assign Brxvx4 = (~(Nxxvx4 ^ N3svx4));
assign Nxxvx4 = (!Ysxvx4);
assign Ysxvx4 = (Gxxvx4 ^ C1svx4);
assign Gxxvx4 = (~(Xvxvx4 ^ Ryrvx4));
assign Xvxvx4 = (Zwxvx4 ^ P39vx4);
assign Zwxvx4 = (Swxvx4 ^ I29vx4);
assign Swxvx4 = (Uz8vx4 ^ B19vx4);
assign Rlxvx4 = (Uxxvx4 & Byxvx4);
assign Byxvx4 = (~(Zpqvx4 & I29vx4));
assign Zpqvx4 = (Ukpvx4 & Iyxvx4);
assign Iyxvx4 = (Pyxvx4 | Lxwvx4);
assign Uxxvx4 = (~(Lrevx4 & Irqvx4));
assign Irqvx4 = (~(Wyxvx4 | Aopvx4));
assign Aopvx4 = (Agxvx4 & Dzxvx4);
assign Dzxvx4 = (~(Kzxvx4 & Gcqvx4));
assign Dlxvx4 = (Rzxvx4 & Yzxvx4);
assign Yzxvx4 = (F0yvx4 & M0yvx4);
assign M0yvx4 = (Uasvx4 | Qaxvx4);
assign Qaxvx4 = (T0yvx4 & A1yvx4);
assign A1yvx4 = (~(H1yvx4 & Lcpvx4));
assign H1yvx4 = (~(O1yvx4 & Ciwvx4));
assign Ciwvx4 = (~(V1yvx4 & C2yvx4));
assign T0yvx4 = (Xaxvx4 | Ud9vx4);
assign F0yvx4 = (~(P39vx4 & Rmpvx4));
assign Rmpvx4 = (~(J2yvx4 & Q2yvx4));
assign Q2yvx4 = (X2yvx4 & E3yvx4);
assign E3yvx4 = (~(L3yvx4 & S3yvx4));
assign S3yvx4 = (~(Qfsvx4 | Aj9vx4));
assign L3yvx4 = (Ukpvx4 & Xhxvx4);
assign X2yvx4 = (~(Ohwvx4 & Fdsvx4));
assign J2yvx4 = (Z3yvx4 & G4yvx4);
assign G4yvx4 = (N4yvx4 | U4yvx4);
assign Rzxvx4 = (B5yvx4 & I5yvx4);
assign I5yvx4 = (~(Dsqvx4 & Y99vx4));
assign B5yvx4 = (~(P5yvx4 & W5yvx4));
assign G2mvx4 = (K6yvx4 ? D6yvx4 : Fs8vx4);
assign D6yvx4 = (~(R6yvx4 & Y6yvx4));
assign Y6yvx4 = (F7yvx4 & M7yvx4);
assign M7yvx4 = (T7yvx4 & A8yvx4);
assign T7yvx4 = (~(H8yvx4 & B19vx4));
assign F7yvx4 = (O8yvx4 & V8yvx4);
assign V8yvx4 = (~(C9yvx4 & J9yvx4));
assign J9yvx4 = (~(Q9yvx4 & X9yvx4));
assign Q9yvx4 = (Sayvx4 ? Layvx4 : Eayvx4);
assign Eayvx4 = (Ot9vx4 | Su9vx4);
assign O8yvx4 = (~(W49vx4 & Zayvx4));
assign R6yvx4 = (Gbyvx4 & Nbyvx4);
assign Gbyvx4 = (Ubyvx4 & Bcyvx4);
assign Bcyvx4 = (Icyvx4 | Y5svx4);
assign Ubyvx4 = (~(Su9vx4 & Pcyvx4));
assign Z1mvx4 = (Wcyvx4 ? J3qvx4 : vis_r2_o[31]);
assign S1mvx4 = (Wcyvx4 ? C3qvx4 : vis_r2_o[28]);
assign L1mvx4 = (Wcyvx4 ? Z4qvx4 : vis_r2_o[7]);
assign E1mvx4 = (Wcyvx4 ? Qppvx4 : vis_r2_o[1]);
assign X0mvx4 = (Wcyvx4 ? G5qvx4 : vis_r2_o[0]);
assign Q0mvx4 = (Ddyvx4 ? J3qvx4 : vis_r3_o[31]);
assign J0mvx4 = (Ddyvx4 ? C3qvx4 : vis_r3_o[28]);
assign C0mvx4 = (Ddyvx4 ? Z4qvx4 : vis_r3_o[7]);
assign Vzlvx4 = (Ddyvx4 ? Qppvx4 : vis_r3_o[1]);
assign Ozlvx4 = (Ddyvx4 ? G5qvx4 : vis_r3_o[0]);
assign Hzlvx4 = (Kdyvx4 ? J3qvx4 : vis_r8_o[31]);
assign Azlvx4 = (Kdyvx4 ? C3qvx4 : vis_r8_o[28]);
assign Tylvx4 = (Kdyvx4 ? Z4qvx4 : vis_r8_o[7]);
assign Mylvx4 = (Kdyvx4 ? Qppvx4 : vis_r8_o[1]);
assign Fylvx4 = (Kdyvx4 ? G5qvx4 : vis_r8_o[0]);
assign Yxlvx4 = (Rdyvx4 ? J3qvx4 : vis_r9_o[31]);
assign Rxlvx4 = (Rdyvx4 ? C3qvx4 : vis_r9_o[28]);
assign Kxlvx4 = (Rdyvx4 ? Z4qvx4 : vis_r9_o[7]);
assign Dxlvx4 = (Rdyvx4 ? Qppvx4 : vis_r9_o[1]);
assign Wwlvx4 = (Rdyvx4 ? G5qvx4 : vis_r9_o[0]);
assign Pwlvx4 = (Ydyvx4 ? J3qvx4 : vis_r10_o[31]);
assign Iwlvx4 = (Ydyvx4 ? C3qvx4 : vis_r10_o[28]);
assign Bwlvx4 = (Ydyvx4 ? Z4qvx4 : vis_r10_o[7]);
assign Uvlvx4 = (Ydyvx4 ? Qppvx4 : vis_r10_o[1]);
assign Nvlvx4 = (Ydyvx4 ? G5qvx4 : vis_r10_o[0]);
assign Gvlvx4 = (Feyvx4 ? J3qvx4 : vis_r11_o[31]);
assign Zulvx4 = (Feyvx4 ? C3qvx4 : vis_r11_o[28]);
assign Sulvx4 = (Feyvx4 ? Z4qvx4 : vis_r11_o[7]);
assign Lulvx4 = (Feyvx4 ? Qppvx4 : vis_r11_o[1]);
assign Eulvx4 = (Feyvx4 ? G5qvx4 : vis_r11_o[0]);
assign Xtlvx4 = (Meyvx4 ? J3qvx4 : vis_r14_o[31]);
assign Qtlvx4 = (Meyvx4 ? C3qvx4 : vis_r14_o[28]);
assign Jtlvx4 = (Meyvx4 ? Z4qvx4 : vis_r14_o[7]);
assign Ctlvx4 = (Meyvx4 ? Qppvx4 : vis_r14_o[1]);
assign Vslvx4 = (Meyvx4 ? G5qvx4 : vis_r14_o[0]);
assign Oslvx4 = (Teyvx4 ? J3qvx4 : vis_r12_o[31]);
assign Hslvx4 = (Teyvx4 ? C3qvx4 : vis_r12_o[28]);
assign Aslvx4 = (Teyvx4 ? Z4qvx4 : vis_r12_o[7]);
assign Trlvx4 = (Teyvx4 ? Qppvx4 : vis_r12_o[1]);
assign Mrlvx4 = (Teyvx4 ? G5qvx4 : vis_r12_o[0]);
assign Frlvx4 = (Afyvx4 ? J3qvx4 : vis_r7_o[31]);
assign Yqlvx4 = (Afyvx4 ? C3qvx4 : vis_r7_o[28]);
assign Rqlvx4 = (Afyvx4 ? Z4qvx4 : vis_r7_o[7]);
assign Kqlvx4 = (Afyvx4 ? Qppvx4 : vis_r7_o[1]);
assign Dqlvx4 = (Afyvx4 ? G5qvx4 : vis_r7_o[0]);
assign Wplvx4 = (Hfyvx4 ? J3qvx4 : vis_r6_o[31]);
assign Pplvx4 = (Hfyvx4 ? C3qvx4 : vis_r6_o[28]);
assign Iplvx4 = (Hfyvx4 ? Z4qvx4 : vis_r6_o[7]);
assign Bplvx4 = (Hfyvx4 ? Qppvx4 : vis_r6_o[1]);
assign Uolvx4 = (Hfyvx4 ? G5qvx4 : vis_r6_o[0]);
assign Nolvx4 = (Ofyvx4 ? J3qvx4 : vis_r5_o[31]);
assign Golvx4 = (Ofyvx4 ? C3qvx4 : vis_r5_o[28]);
assign Znlvx4 = (Ofyvx4 ? Z4qvx4 : vis_r5_o[7]);
assign Snlvx4 = (Ofyvx4 ? Qppvx4 : vis_r5_o[1]);
assign Lnlvx4 = (Ofyvx4 ? G5qvx4 : vis_r5_o[0]);
assign Enlvx4 = (Vfyvx4 ? J3qvx4 : vis_r4_o[31]);
assign Xmlvx4 = (Vfyvx4 ? C3qvx4 : vis_r4_o[28]);
assign Qmlvx4 = (Vfyvx4 ? Z4qvx4 : vis_r4_o[7]);
assign Jmlvx4 = (Vfyvx4 ? Qppvx4 : vis_r4_o[1]);
assign Qppvx4 = (~(C2rvx4 & Cgyvx4));
assign Cmlvx4 = (Vfyvx4 ? G5qvx4 : vis_r4_o[0]);
assign G5qvx4 = (~(Jgyvx4 & Qgyvx4));
assign Qgyvx4 = (Xgyvx4 & Ehyvx4);
assign Ehyvx4 = (~(Dmh2z4[0] & Lhyvx4));
assign Xgyvx4 = (Shyvx4 | Zhyvx4);
assign Jgyvx4 = (~(Giyvx4 | F9pvx4));
assign F9pvx4 = (~(Niyvx4 & Uiyvx4));
assign Uiyvx4 = (Bjyvx4 & Ijyvx4);
assign Ijyvx4 = (~(Pjyvx4 & Wjyvx4));
assign Bjyvx4 = (Dkyvx4 & Kkyvx4);
assign Dkyvx4 = (~(Rkyvx4 & Ykyvx4));
assign Niyvx4 = (Flyvx4 & Mlyvx4);
assign Mlyvx4 = (~(Tlyvx4 & Amyvx4));
assign Flyvx4 = (~(Hmyvx4 & Omyvx4));
assign Vllvx4 = (~(Vmyvx4 & Cnyvx4));
assign Cnyvx4 = (Jnyvx4 & Qnyvx4);
assign Qnyvx4 = (~(Xnyvx4 & Eoyvx4));
assign Eoyvx4 = (~(Loyvx4 | Soyvx4));
assign Xnyvx4 = (~(R1pvx4 | Qoxvx4));
assign Jnyvx4 = (~(P0pvx4 & vis_ipsr_o[1]));
assign Vmyvx4 = (Zoyvx4 & Gpyvx4);
assign Gpyvx4 = (~(W0pvx4 & vis_pc_o[0]));
assign Zoyvx4 = (~(Uzcvx4 & F2pvx4));
assign Ollvx4 = (Upyvx4 ? Npyvx4 : vis_control_o);
assign Upyvx4 = (Bqyvx4 & hready_i);
assign Bqyvx4 = (~(Iqyvx4 & Pqyvx4));
assign Pqyvx4 = (~(Wqyvx4 & Dryvx4));
assign Dryvx4 = (Yo9vx4 & Kryvx4);
assign Wqyvx4 = (~(Rryvx4 | Yryvx4));
assign Iqyvx4 = (~(Fsyvx4 | Msyvx4));
assign Npyvx4 = (~(Tsyvx4 & Atyvx4));
assign Atyvx4 = (~(Kryvx4 & Htyvx4));
assign Tsyvx4 = (~(Hx8vx4 & vis_pc_o[1]));
assign Hllvx4 = (Vtyvx4 ? Otyvx4 : O7evx4);
assign Vtyvx4 = (Cuyvx4 & hready_i);
assign Cuyvx4 = (~(Juyvx4 & Quyvx4));
assign Quyvx4 = (Xuyvx4 & Evyvx4);
assign Evyvx4 = (Lvyvx4 & Svyvx4);
assign Lvyvx4 = (Zvyvx4 & Gwyvx4);
assign Xuyvx4 = (Nwyvx4 & Uwyvx4);
assign Uwyvx4 = (~(Bxyvx4 & Ffqvx4));
assign Nwyvx4 = (~(Ixyvx4 & Wdqvx4));
assign Ixyvx4 = (~(Pxyvx4 | Vdgvx4));
assign Juyvx4 = (Wxyvx4 & Dyyvx4);
assign Dyyvx4 = (Kyyvx4 & Ryyvx4);
assign Ryyvx4 = (Yyyvx4 | Fjgvx4);
assign Kyyvx4 = (Fzyvx4 | Gwrvx4);
assign Wxyvx4 = (Mzyvx4 & Tzyvx4);
assign Tzyvx4 = (~(P5yvx4 & Eznvx4));
assign Mzyvx4 = (~(A0zvx4 & H0zvx4));
assign Otyvx4 = (~(O0zvx4 & V0zvx4));
assign V0zvx4 = (~(C1zvx4 & J1zvx4));
assign J1zvx4 = (Q1zvx4 | X1zvx4);
assign X1zvx4 = (M3ovx4 ? P6xvx4 : E2zvx4);
assign E2zvx4 = (~(Uz8vx4 & Fjgvx4));
assign Q1zvx4 = (~(L2zvx4 & Bswvx4));
assign L2zvx4 = (Z6gvx4 ? Efgvx4 : P39vx4);
assign C1zvx4 = (vis_control_o | S2zvx4);
assign S2zvx4 = (~(Z2zvx4 | Pnnvx4));
assign O0zvx4 = (Uz8vx4 ? N3zvx4 : G3zvx4);
assign N3zvx4 = (U4yvx4 | Mcgvx4);
assign G3zvx4 = (~(U3zvx4 & B4zvx4));
assign U3zvx4 = (B19vx4 & P39vx4);
assign Allvx4 = (I4zvx4 ? Z4qvx4 : vis_psp_o[5]);
assign Tklvx4 = (I4zvx4 ? C3qvx4 : vis_psp_o[26]);
assign Mklvx4 = (I4zvx4 ? J3qvx4 : vis_psp_o[29]);
assign Fklvx4 = (P4zvx4 ? Z4qvx4 : vis_msp_o[5]);
assign Z4qvx4 = (W4zvx4 | D5zvx4);
assign Yjlvx4 = (P4zvx4 ? C3qvx4 : vis_msp_o[26]);
assign C3qvx4 = (~(K5zvx4 & Wzpvx4));
assign Rjlvx4 = (P4zvx4 ? J3qvx4 : vis_msp_o[29]);
assign J3qvx4 = (~(R5zvx4 & Y5zvx4));
assign Kjlvx4 = (I4zvx4 ? F6zvx4 : vis_psp_o[28]);
assign Djlvx4 = (P4zvx4 ? F6zvx4 : vis_msp_o[28]);
assign Wilvx4 = (Meyvx4 ? F6zvx4 : vis_r14_o[30]);
assign Pilvx4 = (Teyvx4 ? F6zvx4 : vis_r12_o[30]);
assign Iilvx4 = (Afyvx4 ? F6zvx4 : vis_r7_o[30]);
assign Bilvx4 = (Hfyvx4 ? F6zvx4 : vis_r6_o[30]);
assign Uhlvx4 = (Ofyvx4 ? F6zvx4 : vis_r5_o[30]);
assign Nhlvx4 = (Vfyvx4 ? F6zvx4 : vis_r4_o[30]);
assign Ghlvx4 = (Feyvx4 ? F6zvx4 : vis_r11_o[30]);
assign Zglvx4 = (Ydyvx4 ? F6zvx4 : vis_r10_o[30]);
assign Sglvx4 = (Rdyvx4 ? F6zvx4 : vis_r9_o[30]);
assign Lglvx4 = (Kdyvx4 ? F6zvx4 : vis_r8_o[30]);
assign Eglvx4 = (Ddyvx4 ? F6zvx4 : vis_r3_o[30]);
assign Xflvx4 = (Wcyvx4 ? F6zvx4 : vis_r2_o[30]);
assign Qflvx4 = (Siqvx4 ? F6zvx4 : vis_r1_o[30]);
assign Jflvx4 = (Xppvx4 ? F6zvx4 : vis_r0_o[30]);
assign F6zvx4 = (~(M6zvx4 & T6zvx4));
assign T6zvx4 = (A7zvx4 & H7zvx4);
assign H7zvx4 = (Shyvx4 | O7zvx4);
assign A7zvx4 = (V7zvx4 & C8zvx4);
assign C8zvx4 = (~(J8zvx4 & Q8zvx4));
assign J8zvx4 = (Dih2z4 & X8zvx4);
assign V7zvx4 = (~(Dmh2z4[30] & Lhyvx4));
assign M6zvx4 = (E9zvx4 & L9zvx4);
assign Cflvx4 = (Z9zvx4 ? vis_apsr_o[2] : S9zvx4);
assign S9zvx4 = (~(Gazvx4 & Nazvx4));
assign Nazvx4 = (X4pvx4 | E9zvx4);
assign Gazvx4 = (Uazvx4 & Bbzvx4);
assign Bbzvx4 = (~(Wspvx4 & Ibzvx4));
assign Uazvx4 = (Ktpvx4 | O7zvx4);
assign Velvx4 = (~(Pbzvx4 & Wbzvx4));
assign Wbzvx4 = (Dczvx4 & Kczvx4);
assign Kczvx4 = (~(vis_apsr_o[2] & P0pvx4));
assign Dczvx4 = (~(W0pvx4 & vis_pc_o[29]));
assign Pbzvx4 = (Rczvx4 & Yczvx4);
assign Yczvx4 = (~(H3wvx4 & haddr_o[30]));
assign Rczvx4 = (~(S4evx4 & F2pvx4));
assign Oelvx4 = (I4zvx4 ? Fdzvx4 : vis_psp_o[27]);
assign Helvx4 = (P4zvx4 ? Fdzvx4 : vis_msp_o[27]);
assign Aelvx4 = (Meyvx4 ? Fdzvx4 : vis_r14_o[29]);
assign Tdlvx4 = (Teyvx4 ? Fdzvx4 : vis_r12_o[29]);
assign Mdlvx4 = (Afyvx4 ? Fdzvx4 : vis_r7_o[29]);
assign Fdlvx4 = (Hfyvx4 ? Fdzvx4 : vis_r6_o[29]);
assign Yclvx4 = (Ofyvx4 ? Fdzvx4 : vis_r5_o[29]);
assign Rclvx4 = (Vfyvx4 ? Fdzvx4 : vis_r4_o[29]);
assign Kclvx4 = (Feyvx4 ? Fdzvx4 : vis_r11_o[29]);
assign Dclvx4 = (Ydyvx4 ? Fdzvx4 : vis_r10_o[29]);
assign Wblvx4 = (Rdyvx4 ? Fdzvx4 : vis_r9_o[29]);
assign Pblvx4 = (Kdyvx4 ? Fdzvx4 : vis_r8_o[29]);
assign Iblvx4 = (Ddyvx4 ? Fdzvx4 : vis_r3_o[29]);
assign Bblvx4 = (Wcyvx4 ? Fdzvx4 : vis_r2_o[29]);
assign Ualvx4 = (Siqvx4 ? Fdzvx4 : vis_r1_o[29]);
assign Nalvx4 = (Xppvx4 ? Fdzvx4 : vis_r0_o[29]);
assign Fdzvx4 = (~(Bspvx4 & Mdzvx4));
assign Galvx4 = (~(Tdzvx4 & Aezvx4));
assign Aezvx4 = (~(L0evx4 & F2pvx4));
assign Tdzvx4 = (Hezvx4 & Oezvx4);
assign Oezvx4 = (~(vis_pc_o[26] & W0pvx4));
assign Hezvx4 = (R1pvx4 | Vezvx4);
assign Z9lvx4 = (I4zvx4 ? Cfzvx4 : vis_psp_o[25]);
assign S9lvx4 = (P4zvx4 ? Cfzvx4 : vis_msp_o[25]);
assign L9lvx4 = (Meyvx4 ? Cfzvx4 : vis_r14_o[27]);
assign E9lvx4 = (Teyvx4 ? Cfzvx4 : vis_r12_o[27]);
assign X8lvx4 = (Afyvx4 ? Cfzvx4 : vis_r7_o[27]);
assign Q8lvx4 = (Hfyvx4 ? Cfzvx4 : vis_r6_o[27]);
assign J8lvx4 = (Ofyvx4 ? Cfzvx4 : vis_r5_o[27]);
assign C8lvx4 = (Vfyvx4 ? Cfzvx4 : vis_r4_o[27]);
assign V7lvx4 = (Feyvx4 ? Cfzvx4 : vis_r11_o[27]);
assign O7lvx4 = (Ydyvx4 ? Cfzvx4 : vis_r10_o[27]);
assign H7lvx4 = (Rdyvx4 ? Cfzvx4 : vis_r9_o[27]);
assign A7lvx4 = (Kdyvx4 ? Cfzvx4 : vis_r8_o[27]);
assign T6lvx4 = (Ddyvx4 ? Cfzvx4 : vis_r3_o[27]);
assign M6lvx4 = (Wcyvx4 ? Cfzvx4 : vis_r2_o[27]);
assign F6lvx4 = (Siqvx4 ? Cfzvx4 : vis_r1_o[27]);
assign Y5lvx4 = (Xppvx4 ? Cfzvx4 : vis_r0_o[27]);
assign Cfzvx4 = (~(Jfzvx4 & Qfzvx4));
assign Jfzvx4 = (Xfzvx4 & Egzvx4);
assign R5lvx4 = (~(Lgzvx4 & Sgzvx4));
assign Sgzvx4 = (~(Azdvx4 & F2pvx4));
assign Lgzvx4 = (Zgzvx4 & Ghzvx4);
assign Ghzvx4 = (~(vis_pc_o[25] & W0pvx4));
assign Zgzvx4 = (R1pvx4 | Nhzvx4);
assign K5lvx4 = (I4zvx4 ? Uhzvx4 : vis_psp_o[24]);
assign D5lvx4 = (P4zvx4 ? Uhzvx4 : vis_msp_o[24]);
assign W4lvx4 = (Meyvx4 ? Uhzvx4 : vis_r14_o[26]);
assign P4lvx4 = (Teyvx4 ? Uhzvx4 : vis_r12_o[26]);
assign I4lvx4 = (Afyvx4 ? Uhzvx4 : vis_r7_o[26]);
assign B4lvx4 = (Hfyvx4 ? Uhzvx4 : vis_r6_o[26]);
assign U3lvx4 = (Ofyvx4 ? Uhzvx4 : vis_r5_o[26]);
assign N3lvx4 = (Vfyvx4 ? Uhzvx4 : vis_r4_o[26]);
assign G3lvx4 = (Feyvx4 ? Uhzvx4 : vis_r11_o[26]);
assign Z2lvx4 = (Ydyvx4 ? Uhzvx4 : vis_r10_o[26]);
assign S2lvx4 = (Rdyvx4 ? Uhzvx4 : vis_r9_o[26]);
assign L2lvx4 = (Kdyvx4 ? Uhzvx4 : vis_r8_o[26]);
assign E2lvx4 = (Ddyvx4 ? Uhzvx4 : vis_r3_o[26]);
assign X1lvx4 = (Wcyvx4 ? Uhzvx4 : vis_r2_o[26]);
assign Q1lvx4 = (Siqvx4 ? Uhzvx4 : vis_r1_o[26]);
assign J1lvx4 = (Xppvx4 ? Uhzvx4 : vis_r0_o[26]);
assign Uhzvx4 = (~(Bizvx4 & Iizvx4));
assign Iizvx4 = (Pizvx4 & Wizvx4);
assign Wizvx4 = (Shyvx4 | Djzvx4);
assign Pizvx4 = (Kjzvx4 & Egzvx4);
assign Kjzvx4 = (~(Dmh2z4[26] & Lhyvx4));
assign Bizvx4 = (Rjzvx4 & Yjzvx4);
assign Rjzvx4 = (Vnbvx4 ? Mkzvx4 : Fkzvx4);
assign Mkzvx4 = (Hlzvx4 ? Alzvx4 : Tkzvx4);
assign Fkzvx4 = (Olzvx4 | Hlzvx4);
assign C1lvx4 = (~(Vlzvx4 & Cmzvx4));
assign Cmzvx4 = (~(Pxdvx4 & F2pvx4));
assign Vlzvx4 = (Jmzvx4 & Qmzvx4);
assign Qmzvx4 = (~(vis_pc_o[24] & W0pvx4));
assign Jmzvx4 = (R1pvx4 | Rnovx4);
assign V0lvx4 = (I4zvx4 ? Xmzvx4 : vis_psp_o[23]);
assign O0lvx4 = (P4zvx4 ? Xmzvx4 : vis_msp_o[23]);
assign H0lvx4 = (Meyvx4 ? Xmzvx4 : vis_r14_o[25]);
assign A0lvx4 = (Teyvx4 ? Xmzvx4 : vis_r12_o[25]);
assign Tzkvx4 = (Afyvx4 ? Xmzvx4 : vis_r7_o[25]);
assign Mzkvx4 = (Hfyvx4 ? Xmzvx4 : vis_r6_o[25]);
assign Fzkvx4 = (Ofyvx4 ? Xmzvx4 : vis_r5_o[25]);
assign Yykvx4 = (Vfyvx4 ? Xmzvx4 : vis_r4_o[25]);
assign Rykvx4 = (Feyvx4 ? Xmzvx4 : vis_r11_o[25]);
assign Kykvx4 = (Ydyvx4 ? Xmzvx4 : vis_r10_o[25]);
assign Dykvx4 = (Rdyvx4 ? Xmzvx4 : vis_r9_o[25]);
assign Wxkvx4 = (Kdyvx4 ? Xmzvx4 : vis_r8_o[25]);
assign Pxkvx4 = (Ddyvx4 ? Xmzvx4 : vis_r3_o[25]);
assign Ixkvx4 = (Wcyvx4 ? Xmzvx4 : vis_r2_o[25]);
assign Bxkvx4 = (Siqvx4 ? Xmzvx4 : vis_r1_o[25]);
assign Uwkvx4 = (Xppvx4 ? Xmzvx4 : vis_r0_o[25]);
assign Xmzvx4 = (~(Enzvx4 & Lnzvx4));
assign Lnzvx4 = (Snzvx4 & Znzvx4);
assign Znzvx4 = (~(Gozvx4 & Nozvx4));
assign Gozvx4 = (X8zvx4 & Kmbvx4);
assign Snzvx4 = (~(Uozvx4 | Bpzvx4));
assign Enzvx4 = (Ipzvx4 & Ppzvx4);
assign Ipzvx4 = (Wpzvx4 & Dqzvx4);
assign Dqzvx4 = (~(Dmh2z4[25] & Lhyvx4));
assign Wpzvx4 = (Shyvx4 | Kqzvx4);
assign Nwkvx4 = (I4zvx4 ? Rqzvx4 : vis_psp_o[22]);
assign Gwkvx4 = (P4zvx4 ? Rqzvx4 : vis_msp_o[22]);
assign Zvkvx4 = (Meyvx4 ? Rqzvx4 : vis_r14_o[24]);
assign Svkvx4 = (Teyvx4 ? Rqzvx4 : vis_r12_o[24]);
assign Lvkvx4 = (Afyvx4 ? Rqzvx4 : vis_r7_o[24]);
assign Evkvx4 = (Hfyvx4 ? Rqzvx4 : vis_r6_o[24]);
assign Xukvx4 = (Ofyvx4 ? Rqzvx4 : vis_r5_o[24]);
assign Qukvx4 = (Vfyvx4 ? Rqzvx4 : vis_r4_o[24]);
assign Jukvx4 = (Feyvx4 ? Rqzvx4 : vis_r11_o[24]);
assign Cukvx4 = (Ydyvx4 ? Rqzvx4 : vis_r10_o[24]);
assign Vtkvx4 = (Rdyvx4 ? Rqzvx4 : vis_r9_o[24]);
assign Otkvx4 = (Kdyvx4 ? Rqzvx4 : vis_r8_o[24]);
assign Htkvx4 = (Ddyvx4 ? Rqzvx4 : vis_r3_o[24]);
assign Atkvx4 = (Wcyvx4 ? Rqzvx4 : vis_r2_o[24]);
assign Tskvx4 = (Siqvx4 ? Rqzvx4 : vis_r1_o[24]);
assign Mskvx4 = (Xppvx4 ? Rqzvx4 : vis_r0_o[24]);
assign Rqzvx4 = (~(O3pvx4 & Yqzvx4));
assign Fskvx4 = (~(Frzvx4 & Mrzvx4));
assign Mrzvx4 = (~(S6dvx4 & F2pvx4));
assign Frzvx4 = (Trzvx4 & Aszvx4);
assign Aszvx4 = (~(vis_pc_o[5] & W0pvx4));
assign Trzvx4 = (R1pvx4 | Hszvx4);
assign Yrkvx4 = (I4zvx4 ? Oszvx4 : vis_psp_o[4]);
assign Rrkvx4 = (P4zvx4 ? Oszvx4 : vis_msp_o[4]);
assign Krkvx4 = (Meyvx4 ? Oszvx4 : vis_r14_o[6]);
assign Drkvx4 = (Teyvx4 ? Oszvx4 : vis_r12_o[6]);
assign Wqkvx4 = (Afyvx4 ? Oszvx4 : vis_r7_o[6]);
assign Pqkvx4 = (Hfyvx4 ? Oszvx4 : vis_r6_o[6]);
assign Iqkvx4 = (Ofyvx4 ? Oszvx4 : vis_r5_o[6]);
assign Bqkvx4 = (Vfyvx4 ? Oszvx4 : vis_r4_o[6]);
assign Upkvx4 = (Feyvx4 ? Oszvx4 : vis_r11_o[6]);
assign Npkvx4 = (Ydyvx4 ? Oszvx4 : vis_r10_o[6]);
assign Gpkvx4 = (Rdyvx4 ? Oszvx4 : vis_r9_o[6]);
assign Zokvx4 = (Kdyvx4 ? Oszvx4 : vis_r8_o[6]);
assign Sokvx4 = (Ddyvx4 ? Oszvx4 : vis_r3_o[6]);
assign Lokvx4 = (Wcyvx4 ? Oszvx4 : vis_r2_o[6]);
assign Eokvx4 = (Siqvx4 ? Oszvx4 : vis_r1_o[6]);
assign Xnkvx4 = (Xppvx4 ? Oszvx4 : vis_r0_o[6]);
assign Oszvx4 = (~(Vszvx4 & Ctzvx4));
assign Ctzvx4 = (Jtzvx4 & Qtzvx4);
assign Qtzvx4 = (~(Xtzvx4 & Euzvx4));
assign Xtzvx4 = (O2bvx4 & X8zvx4);
assign Jtzvx4 = (Luzvx4 & Egzvx4);
assign Vszvx4 = (Suzvx4 & Zuzvx4);
assign Suzvx4 = (Gvzvx4 & Nvzvx4);
assign Nvzvx4 = (~(Dmh2z4[6] & Lhyvx4));
assign Gvzvx4 = (Shyvx4 | Uvzvx4);
assign Qnkvx4 = (~(Bwzvx4 & Iwzvx4));
assign Iwzvx4 = (Pwzvx4 & Wwzvx4);
assign Wwzvx4 = (~(vis_ipsr_o[5] & P0pvx4));
assign Pwzvx4 = (~(vis_pc_o[4] & W0pvx4));
assign Bwzvx4 = (Dxzvx4 & Kxzvx4);
assign Kxzvx4 = (R1pvx4 | Rxzvx4);
assign Dxzvx4 = (~(I5dvx4 & F2pvx4));
assign Jnkvx4 = (I4zvx4 ? Yxzvx4 : vis_psp_o[3]);
assign Cnkvx4 = (P4zvx4 ? Yxzvx4 : vis_msp_o[3]);
assign Vmkvx4 = (Meyvx4 ? Yxzvx4 : vis_r14_o[5]);
assign Omkvx4 = (Teyvx4 ? Yxzvx4 : vis_r12_o[5]);
assign Hmkvx4 = (Afyvx4 ? Yxzvx4 : vis_r7_o[5]);
assign Amkvx4 = (Hfyvx4 ? Yxzvx4 : vis_r6_o[5]);
assign Tlkvx4 = (Ofyvx4 ? Yxzvx4 : vis_r5_o[5]);
assign Mlkvx4 = (Vfyvx4 ? Yxzvx4 : vis_r4_o[5]);
assign Flkvx4 = (Feyvx4 ? Yxzvx4 : vis_r11_o[5]);
assign Ykkvx4 = (Ydyvx4 ? Yxzvx4 : vis_r10_o[5]);
assign Rkkvx4 = (Rdyvx4 ? Yxzvx4 : vis_r9_o[5]);
assign Kkkvx4 = (Kdyvx4 ? Yxzvx4 : vis_r8_o[5]);
assign Dkkvx4 = (Ddyvx4 ? Yxzvx4 : vis_r3_o[5]);
assign Wjkvx4 = (Wcyvx4 ? Yxzvx4 : vis_r2_o[5]);
assign Pjkvx4 = (Siqvx4 ? Yxzvx4 : vis_r1_o[5]);
assign Ijkvx4 = (Xppvx4 ? Yxzvx4 : vis_r0_o[5]);
assign Yxzvx4 = (~(Vcuvx4 & Fyzvx4));
assign Bjkvx4 = (~(Myzvx4 & Tyzvx4));
assign Tyzvx4 = (Azzvx4 & Hzzvx4);
assign Hzzvx4 = (~(P0pvx4 & vis_ipsr_o[4]));
assign Azzvx4 = (~(vis_pc_o[3] & W0pvx4));
assign Myzvx4 = (Ozzvx4 & Vzzvx4);
assign Vzzvx4 = (R1pvx4 | Yuovx4);
assign Ozzvx4 = (~(Y3dvx4 & F2pvx4));
assign Uikvx4 = (I4zvx4 ? C00wx4 : vis_psp_o[2]);
assign Nikvx4 = (P4zvx4 ? C00wx4 : vis_msp_o[2]);
assign Gikvx4 = (Meyvx4 ? C00wx4 : vis_r14_o[4]);
assign Zhkvx4 = (Teyvx4 ? C00wx4 : vis_r12_o[4]);
assign Shkvx4 = (Afyvx4 ? C00wx4 : vis_r7_o[4]);
assign Lhkvx4 = (Hfyvx4 ? C00wx4 : vis_r6_o[4]);
assign Ehkvx4 = (Ofyvx4 ? C00wx4 : vis_r5_o[4]);
assign Xgkvx4 = (Vfyvx4 ? C00wx4 : vis_r4_o[4]);
assign Qgkvx4 = (Feyvx4 ? C00wx4 : vis_r11_o[4]);
assign Jgkvx4 = (Ydyvx4 ? C00wx4 : vis_r10_o[4]);
assign Cgkvx4 = (Rdyvx4 ? C00wx4 : vis_r9_o[4]);
assign Vfkvx4 = (Kdyvx4 ? C00wx4 : vis_r8_o[4]);
assign Ofkvx4 = (Ddyvx4 ? C00wx4 : vis_r3_o[4]);
assign Hfkvx4 = (Wcyvx4 ? C00wx4 : vis_r2_o[4]);
assign Afkvx4 = (Siqvx4 ? C00wx4 : vis_r1_o[4]);
assign Tekvx4 = (Xppvx4 ? C00wx4 : vis_r0_o[4]);
assign C00wx4 = (~(Leuvx4 & J00wx4));
assign Mekvx4 = (~(Q00wx4 & X00wx4));
assign X00wx4 = (E10wx4 & L10wx4);
assign L10wx4 = (R1pvx4 | Ekovx4);
assign Ekovx4 = (S10wx4 & Z10wx4);
assign Z10wx4 = (~(Gzvvx4 & Aqnvx4));
assign S10wx4 = (G20wx4 & N20wx4);
assign N20wx4 = (~(Ykh2z4[2] & Mrsvx4));
assign G20wx4 = (~(Dmh2z4[3] & K1wvx4));
assign E10wx4 = (~(P0pvx4 & vis_ipsr_o[3]));
assign Q00wx4 = (U20wx4 & B30wx4);
assign B30wx4 = (~(W0pvx4 & vis_pc_o[2]));
assign U20wx4 = (~(O2dvx4 & F2pvx4));
assign Fekvx4 = (I4zvx4 ? I30wx4 : vis_psp_o[1]);
assign Ydkvx4 = (P4zvx4 ? I30wx4 : vis_msp_o[1]);
assign Rdkvx4 = (Meyvx4 ? I30wx4 : vis_r14_o[3]);
assign Kdkvx4 = (Teyvx4 ? I30wx4 : vis_r12_o[3]);
assign Ddkvx4 = (Afyvx4 ? I30wx4 : vis_r7_o[3]);
assign Wckvx4 = (Hfyvx4 ? I30wx4 : vis_r6_o[3]);
assign Pckvx4 = (Ofyvx4 ? I30wx4 : vis_r5_o[3]);
assign Ickvx4 = (Vfyvx4 ? I30wx4 : vis_r4_o[3]);
assign Bckvx4 = (Feyvx4 ? I30wx4 : vis_r11_o[3]);
assign Ubkvx4 = (Ydyvx4 ? I30wx4 : vis_r10_o[3]);
assign Nbkvx4 = (Rdyvx4 ? I30wx4 : vis_r9_o[3]);
assign Gbkvx4 = (Kdyvx4 ? I30wx4 : vis_r8_o[3]);
assign Zakvx4 = (Ddyvx4 ? I30wx4 : vis_r3_o[3]);
assign Sakvx4 = (Wcyvx4 ? I30wx4 : vis_r2_o[3]);
assign Lakvx4 = (Siqvx4 ? I30wx4 : vis_r1_o[3]);
assign Eakvx4 = (Xppvx4 ? I30wx4 : vis_r0_o[3]);
assign I30wx4 = (~(P30wx4 & W30wx4));
assign W30wx4 = (D40wx4 & K40wx4);
assign K40wx4 = (Shyvx4 | R40wx4);
assign D40wx4 = (Y40wx4 & F50wx4);
assign F50wx4 = (Egzvx4 | Rryvx4);
assign Y40wx4 = (~(Dmh2z4[3] & Lhyvx4));
assign P30wx4 = (U0vvx4 & M50wx4);
assign X9kvx4 = (U5qvx4 ? T50wx4 : Zph2z4[1]);
assign U5qvx4 = (hready_i & hprot_o[0]);
assign Q9kvx4 = (~(A60wx4 & H60wx4));
assign H60wx4 = (~(Itdvx4 & F2pvx4));
assign A60wx4 = (O60wx4 & V60wx4);
assign V60wx4 = (~(vis_pc_o[21] & W0pvx4));
assign O60wx4 = (R1pvx4 | C70wx4);
assign J9kvx4 = (I4zvx4 ? J70wx4 : vis_psp_o[20]);
assign C9kvx4 = (P4zvx4 ? J70wx4 : vis_msp_o[20]);
assign V8kvx4 = (Meyvx4 ? J70wx4 : vis_r14_o[22]);
assign O8kvx4 = (Teyvx4 ? J70wx4 : vis_r12_o[22]);
assign H8kvx4 = (Afyvx4 ? J70wx4 : vis_r7_o[22]);
assign A8kvx4 = (Hfyvx4 ? J70wx4 : vis_r6_o[22]);
assign T7kvx4 = (Ofyvx4 ? J70wx4 : vis_r5_o[22]);
assign M7kvx4 = (Vfyvx4 ? J70wx4 : vis_r4_o[22]);
assign F7kvx4 = (Feyvx4 ? J70wx4 : vis_r11_o[22]);
assign Y6kvx4 = (Ydyvx4 ? J70wx4 : vis_r10_o[22]);
assign R6kvx4 = (Rdyvx4 ? J70wx4 : vis_r9_o[22]);
assign K6kvx4 = (Kdyvx4 ? J70wx4 : vis_r8_o[22]);
assign D6kvx4 = (Ddyvx4 ? J70wx4 : vis_r3_o[22]);
assign W5kvx4 = (Wcyvx4 ? J70wx4 : vis_r2_o[22]);
assign P5kvx4 = (Siqvx4 ? J70wx4 : vis_r1_o[22]);
assign I5kvx4 = (Xppvx4 ? J70wx4 : vis_r0_o[22]);
assign J70wx4 = (~(Q70wx4 & X70wx4));
assign X70wx4 = (E80wx4 & L80wx4);
assign L80wx4 = (~(Dmh2z4[22] & Lhyvx4));
assign E80wx4 = (S80wx4 & Z80wx4);
assign S80wx4 = (~(G90wx4 & N90wx4));
assign G90wx4 = (Zkbvx4 & X8zvx4);
assign Q70wx4 = (U90wx4 & Ba0wx4);
assign U90wx4 = (Ia0wx4 & Pa0wx4);
assign Pa0wx4 = (Shyvx4 | Wa0wx4);
assign B5kvx4 = (~(Db0wx4 & Kb0wx4));
assign Kb0wx4 = (~(Xrdvx4 & F2pvx4));
assign Db0wx4 = (Rb0wx4 & Yb0wx4);
assign Yb0wx4 = (~(vis_pc_o[20] & W0pvx4));
assign Rb0wx4 = (R1pvx4 | Fc0wx4);
assign U4kvx4 = (I4zvx4 ? Mc0wx4 : vis_psp_o[19]);
assign N4kvx4 = (P4zvx4 ? Mc0wx4 : vis_msp_o[19]);
assign G4kvx4 = (Meyvx4 ? Mc0wx4 : vis_r14_o[21]);
assign Z3kvx4 = (Teyvx4 ? Mc0wx4 : vis_r12_o[21]);
assign S3kvx4 = (Afyvx4 ? Mc0wx4 : vis_r7_o[21]);
assign L3kvx4 = (Hfyvx4 ? Mc0wx4 : vis_r6_o[21]);
assign E3kvx4 = (Ofyvx4 ? Mc0wx4 : vis_r5_o[21]);
assign X2kvx4 = (Vfyvx4 ? Mc0wx4 : vis_r4_o[21]);
assign Q2kvx4 = (Feyvx4 ? Mc0wx4 : vis_r11_o[21]);
assign J2kvx4 = (Ydyvx4 ? Mc0wx4 : vis_r10_o[21]);
assign C2kvx4 = (Rdyvx4 ? Mc0wx4 : vis_r9_o[21]);
assign V1kvx4 = (Kdyvx4 ? Mc0wx4 : vis_r8_o[21]);
assign O1kvx4 = (Ddyvx4 ? Mc0wx4 : vis_r3_o[21]);
assign H1kvx4 = (Wcyvx4 ? Mc0wx4 : vis_r2_o[21]);
assign A1kvx4 = (Siqvx4 ? Mc0wx4 : vis_r1_o[21]);
assign T0kvx4 = (Xppvx4 ? Mc0wx4 : vis_r0_o[21]);
assign Mc0wx4 = (~(Tc0wx4 & Ad0wx4));
assign Ad0wx4 = (Hd0wx4 & Ia0wx4);
assign Hd0wx4 = (Od0wx4 & Vd0wx4);
assign Vd0wx4 = (~(Dmh2z4[21] & Lhyvx4));
assign Od0wx4 = (Shyvx4 | Ce0wx4);
assign Tc0wx4 = (Je0wx4 & Qe0wx4);
assign Je0wx4 = (Ojbvx4 ? Ef0wx4 : Xe0wx4);
assign Ef0wx4 = (Lf0wx4 ? Alzvx4 : Tkzvx4);
assign Xe0wx4 = (Olzvx4 | Lf0wx4);
assign M0kvx4 = (~(Sf0wx4 & Zf0wx4));
assign Zf0wx4 = (~(Mqdvx4 & F2pvx4));
assign Sf0wx4 = (Gg0wx4 & Ng0wx4);
assign Ng0wx4 = (~(vis_pc_o[19] & W0pvx4));
assign Gg0wx4 = (R1pvx4 | Ug0wx4);
assign F0kvx4 = (I4zvx4 ? Bh0wx4 : vis_psp_o[18]);
assign Yzjvx4 = (P4zvx4 ? Bh0wx4 : vis_msp_o[18]);
assign Rzjvx4 = (Meyvx4 ? Bh0wx4 : vis_r14_o[20]);
assign Kzjvx4 = (Teyvx4 ? Bh0wx4 : vis_r12_o[20]);
assign Dzjvx4 = (Afyvx4 ? Bh0wx4 : vis_r7_o[20]);
assign Wyjvx4 = (Hfyvx4 ? Bh0wx4 : vis_r6_o[20]);
assign Pyjvx4 = (Ofyvx4 ? Bh0wx4 : vis_r5_o[20]);
assign Iyjvx4 = (Vfyvx4 ? Bh0wx4 : vis_r4_o[20]);
assign Byjvx4 = (Feyvx4 ? Bh0wx4 : vis_r11_o[20]);
assign Uxjvx4 = (Ydyvx4 ? Bh0wx4 : vis_r10_o[20]);
assign Nxjvx4 = (Rdyvx4 ? Bh0wx4 : vis_r9_o[20]);
assign Gxjvx4 = (Kdyvx4 ? Bh0wx4 : vis_r8_o[20]);
assign Zwjvx4 = (Ddyvx4 ? Bh0wx4 : vis_r3_o[20]);
assign Swjvx4 = (Wcyvx4 ? Bh0wx4 : vis_r2_o[20]);
assign Lwjvx4 = (Siqvx4 ? Bh0wx4 : vis_r1_o[20]);
assign Ewjvx4 = (Xppvx4 ? Bh0wx4 : vis_r0_o[20]);
assign Bh0wx4 = (~(Ih0wx4 & Ph0wx4));
assign Ph0wx4 = (Wh0wx4 & Di0wx4);
assign Di0wx4 = (~(Dmh2z4[20] & Lhyvx4));
assign Wh0wx4 = (Ki0wx4 & Ri0wx4);
assign Ki0wx4 = (~(Yi0wx4 & Fj0wx4));
assign Yi0wx4 = (Dibvx4 & X8zvx4);
assign Ih0wx4 = (Mj0wx4 & Tj0wx4);
assign Mj0wx4 = (Ia0wx4 & Ak0wx4);
assign Ak0wx4 = (Shyvx4 | Hk0wx4);
assign Xvjvx4 = (~(Ok0wx4 & Vk0wx4));
assign Vk0wx4 = (~(Bpdvx4 & F2pvx4));
assign Ok0wx4 = (Cl0wx4 & Jl0wx4);
assign Jl0wx4 = (~(vis_pc_o[18] & W0pvx4));
assign Cl0wx4 = (R1pvx4 | Ql0wx4);
assign Qvjvx4 = (I4zvx4 ? Xl0wx4 : vis_psp_o[17]);
assign Jvjvx4 = (P4zvx4 ? Xl0wx4 : vis_msp_o[17]);
assign Cvjvx4 = (Meyvx4 ? Xl0wx4 : vis_r14_o[19]);
assign Vujvx4 = (Teyvx4 ? Xl0wx4 : vis_r12_o[19]);
assign Oujvx4 = (Afyvx4 ? Xl0wx4 : vis_r7_o[19]);
assign Hujvx4 = (Hfyvx4 ? Xl0wx4 : vis_r6_o[19]);
assign Aujvx4 = (Ofyvx4 ? Xl0wx4 : vis_r5_o[19]);
assign Ttjvx4 = (Vfyvx4 ? Xl0wx4 : vis_r4_o[19]);
assign Mtjvx4 = (Feyvx4 ? Xl0wx4 : vis_r11_o[19]);
assign Ftjvx4 = (Ydyvx4 ? Xl0wx4 : vis_r10_o[19]);
assign Ysjvx4 = (Rdyvx4 ? Xl0wx4 : vis_r9_o[19]);
assign Rsjvx4 = (Kdyvx4 ? Xl0wx4 : vis_r8_o[19]);
assign Ksjvx4 = (Ddyvx4 ? Xl0wx4 : vis_r3_o[19]);
assign Dsjvx4 = (Wcyvx4 ? Xl0wx4 : vis_r2_o[19]);
assign Wrjvx4 = (Siqvx4 ? Xl0wx4 : vis_r1_o[19]);
assign Prjvx4 = (Xppvx4 ? Xl0wx4 : vis_r0_o[19]);
assign Xl0wx4 = (~(Em0wx4 & Lm0wx4));
assign Lm0wx4 = (Sm0wx4 & Ia0wx4);
assign Sm0wx4 = (Zm0wx4 & Gn0wx4);
assign Gn0wx4 = (~(Dmh2z4[19] & Lhyvx4));
assign Zm0wx4 = (Shyvx4 | Nn0wx4);
assign Em0wx4 = (Un0wx4 & Bo0wx4);
assign Un0wx4 = (Sgbvx4 ? Po0wx4 : Io0wx4);
assign Po0wx4 = (Wo0wx4 ? Alzvx4 : Tkzvx4);
assign Io0wx4 = (Olzvx4 | Wo0wx4);
assign Irjvx4 = (~(Dp0wx4 & Kp0wx4));
assign Kp0wx4 = (~(Qndvx4 & F2pvx4));
assign Dp0wx4 = (Rp0wx4 & Yp0wx4);
assign Yp0wx4 = (~(vis_pc_o[17] & W0pvx4));
assign Rp0wx4 = (R1pvx4 | Fq0wx4);
assign Brjvx4 = (I4zvx4 ? Mq0wx4 : vis_psp_o[16]);
assign Uqjvx4 = (P4zvx4 ? Mq0wx4 : vis_msp_o[16]);
assign Nqjvx4 = (Meyvx4 ? Mq0wx4 : vis_r14_o[18]);
assign Gqjvx4 = (Teyvx4 ? Mq0wx4 : vis_r12_o[18]);
assign Zpjvx4 = (Afyvx4 ? Mq0wx4 : vis_r7_o[18]);
assign Spjvx4 = (Hfyvx4 ? Mq0wx4 : vis_r6_o[18]);
assign Lpjvx4 = (Ofyvx4 ? Mq0wx4 : vis_r5_o[18]);
assign Epjvx4 = (Vfyvx4 ? Mq0wx4 : vis_r4_o[18]);
assign Xojvx4 = (Feyvx4 ? Mq0wx4 : vis_r11_o[18]);
assign Qojvx4 = (Ydyvx4 ? Mq0wx4 : vis_r10_o[18]);
assign Jojvx4 = (Rdyvx4 ? Mq0wx4 : vis_r9_o[18]);
assign Cojvx4 = (Kdyvx4 ? Mq0wx4 : vis_r8_o[18]);
assign Vnjvx4 = (Ddyvx4 ? Mq0wx4 : vis_r3_o[18]);
assign Onjvx4 = (Wcyvx4 ? Mq0wx4 : vis_r2_o[18]);
assign Hnjvx4 = (Siqvx4 ? Mq0wx4 : vis_r1_o[18]);
assign Anjvx4 = (Xppvx4 ? Mq0wx4 : vis_r0_o[18]);
assign Mq0wx4 = (~(Tq0wx4 & Ar0wx4));
assign Ar0wx4 = (Hr0wx4 & Or0wx4);
assign Or0wx4 = (~(Dmh2z4[18] & Lhyvx4));
assign Hr0wx4 = (Vr0wx4 & Cs0wx4);
assign Vr0wx4 = (~(Js0wx4 & Qs0wx4));
assign Js0wx4 = (Hfbvx4 & X8zvx4);
assign Tq0wx4 = (Xs0wx4 & Et0wx4);
assign Xs0wx4 = (Ia0wx4 & Lt0wx4);
assign Lt0wx4 = (Shyvx4 | St0wx4);
assign Tmjvx4 = (~(Zt0wx4 & Gu0wx4));
assign Gu0wx4 = (~(Fmdvx4 & F2pvx4));
assign Zt0wx4 = (Nu0wx4 & Uu0wx4);
assign Uu0wx4 = (~(vis_pc_o[16] & W0pvx4));
assign Nu0wx4 = (R1pvx4 | Bv0wx4);
assign Mmjvx4 = (I4zvx4 ? Iv0wx4 : vis_psp_o[15]);
assign Fmjvx4 = (P4zvx4 ? Iv0wx4 : vis_msp_o[15]);
assign Yljvx4 = (Meyvx4 ? Iv0wx4 : vis_r14_o[17]);
assign Rljvx4 = (Teyvx4 ? Iv0wx4 : vis_r12_o[17]);
assign Kljvx4 = (Afyvx4 ? Iv0wx4 : vis_r7_o[17]);
assign Dljvx4 = (Hfyvx4 ? Iv0wx4 : vis_r6_o[17]);
assign Wkjvx4 = (Ofyvx4 ? Iv0wx4 : vis_r5_o[17]);
assign Pkjvx4 = (Vfyvx4 ? Iv0wx4 : vis_r4_o[17]);
assign Ikjvx4 = (Feyvx4 ? Iv0wx4 : vis_r11_o[17]);
assign Bkjvx4 = (Ydyvx4 ? Iv0wx4 : vis_r10_o[17]);
assign Ujjvx4 = (Rdyvx4 ? Iv0wx4 : vis_r9_o[17]);
assign Njjvx4 = (Kdyvx4 ? Iv0wx4 : vis_r8_o[17]);
assign Gjjvx4 = (Ddyvx4 ? Iv0wx4 : vis_r3_o[17]);
assign Zijvx4 = (Wcyvx4 ? Iv0wx4 : vis_r2_o[17]);
assign Sijvx4 = (Siqvx4 ? Iv0wx4 : vis_r1_o[17]);
assign Lijvx4 = (Xppvx4 ? Iv0wx4 : vis_r0_o[17]);
assign Iv0wx4 = (~(Pv0wx4 & Wv0wx4));
assign Wv0wx4 = (Dw0wx4 & Ia0wx4);
assign Dw0wx4 = (Kw0wx4 & Rw0wx4);
assign Rw0wx4 = (~(Dmh2z4[17] & Lhyvx4));
assign Kw0wx4 = (Shyvx4 | Yw0wx4);
assign Pv0wx4 = (Fx0wx4 & Mx0wx4);
assign Fx0wx4 = (Wdbvx4 ? Ay0wx4 : Tx0wx4);
assign Ay0wx4 = (Hy0wx4 ? Alzvx4 : Tkzvx4);
assign Tx0wx4 = (Olzvx4 | Hy0wx4);
assign Eijvx4 = (~(Oy0wx4 & Vy0wx4));
assign Vy0wx4 = (~(Ukdvx4 & F2pvx4));
assign Oy0wx4 = (Cz0wx4 & Jz0wx4);
assign Jz0wx4 = (~(vis_pc_o[15] & W0pvx4));
assign Cz0wx4 = (R1pvx4 | Vpovx4);
assign Xhjvx4 = (I4zvx4 ? Qz0wx4 : vis_psp_o[14]);
assign Qhjvx4 = (P4zvx4 ? Qz0wx4 : vis_msp_o[14]);
assign Jhjvx4 = (Meyvx4 ? Qz0wx4 : vis_r14_o[16]);
assign Chjvx4 = (Teyvx4 ? Qz0wx4 : vis_r12_o[16]);
assign Vgjvx4 = (Afyvx4 ? Qz0wx4 : vis_r7_o[16]);
assign Ogjvx4 = (Hfyvx4 ? Qz0wx4 : vis_r6_o[16]);
assign Hgjvx4 = (Ofyvx4 ? Qz0wx4 : vis_r5_o[16]);
assign Agjvx4 = (Vfyvx4 ? Qz0wx4 : vis_r4_o[16]);
assign Tfjvx4 = (Feyvx4 ? Qz0wx4 : vis_r11_o[16]);
assign Mfjvx4 = (Ydyvx4 ? Qz0wx4 : vis_r10_o[16]);
assign Ffjvx4 = (Rdyvx4 ? Qz0wx4 : vis_r9_o[16]);
assign Yejvx4 = (Kdyvx4 ? Qz0wx4 : vis_r8_o[16]);
assign Rejvx4 = (Ddyvx4 ? Qz0wx4 : vis_r3_o[16]);
assign Kejvx4 = (Wcyvx4 ? Qz0wx4 : vis_r2_o[16]);
assign Dejvx4 = (Siqvx4 ? Qz0wx4 : vis_r1_o[16]);
assign Wdjvx4 = (Xppvx4 ? Qz0wx4 : vis_r0_o[16]);
assign Qz0wx4 = (~(Xz0wx4 & E01wx4));
assign E01wx4 = (L01wx4 & S01wx4);
assign S01wx4 = (~(Dmh2z4[16] & Lhyvx4));
assign L01wx4 = (Z01wx4 & G11wx4);
assign Z01wx4 = (~(N11wx4 & U11wx4));
assign N11wx4 = (Lcbvx4 & X8zvx4);
assign Xz0wx4 = (B21wx4 & I21wx4);
assign B21wx4 = (Ia0wx4 & P21wx4);
assign P21wx4 = (Shyvx4 | W21wx4);
assign Ia0wx4 = (D31wx4 & Egzvx4);
assign Pdjvx4 = (~(K31wx4 & R31wx4));
assign R31wx4 = (~(Yhdvx4 & F2pvx4));
assign K31wx4 = (Y31wx4 & F41wx4);
assign F41wx4 = (~(vis_pc_o[13] & W0pvx4));
assign Y31wx4 = (~(H3wvx4 & haddr_o[14]));
assign Idjvx4 = (I4zvx4 ? M41wx4 : vis_psp_o[12]);
assign Bdjvx4 = (P4zvx4 ? M41wx4 : vis_msp_o[12]);
assign Ucjvx4 = (Meyvx4 ? M41wx4 : vis_r14_o[14]);
assign Ncjvx4 = (Teyvx4 ? M41wx4 : vis_r12_o[14]);
assign Gcjvx4 = (Afyvx4 ? M41wx4 : vis_r7_o[14]);
assign Zbjvx4 = (Hfyvx4 ? M41wx4 : vis_r6_o[14]);
assign Sbjvx4 = (Ofyvx4 ? M41wx4 : vis_r5_o[14]);
assign Lbjvx4 = (Vfyvx4 ? M41wx4 : vis_r4_o[14]);
assign Ebjvx4 = (Feyvx4 ? M41wx4 : vis_r11_o[14]);
assign Xajvx4 = (Ydyvx4 ? M41wx4 : vis_r10_o[14]);
assign Qajvx4 = (Rdyvx4 ? M41wx4 : vis_r9_o[14]);
assign Jajvx4 = (Kdyvx4 ? M41wx4 : vis_r8_o[14]);
assign Cajvx4 = (Ddyvx4 ? M41wx4 : vis_r3_o[14]);
assign V9jvx4 = (Wcyvx4 ? M41wx4 : vis_r2_o[14]);
assign O9jvx4 = (Siqvx4 ? M41wx4 : vis_r1_o[14]);
assign H9jvx4 = (Xppvx4 ? M41wx4 : vis_r0_o[14]);
assign M41wx4 = (~(T41wx4 & A51wx4));
assign A51wx4 = (H51wx4 & O51wx4);
assign O51wx4 = (~(V51wx4 & C61wx4));
assign V51wx4 = (P9bvx4 & X8zvx4);
assign H51wx4 = (~(J61wx4 | Bpzvx4));
assign T41wx4 = (Q61wx4 & X61wx4);
assign Q61wx4 = (E71wx4 & L71wx4);
assign L71wx4 = (~(Dmh2z4[14] & Lhyvx4));
assign E71wx4 = (Shyvx4 | S71wx4);
assign A9jvx4 = (~(Z71wx4 & G81wx4));
assign G81wx4 = (~(Ngdvx4 & F2pvx4));
assign Z71wx4 = (N81wx4 & U81wx4);
assign U81wx4 = (~(vis_pc_o[12] & W0pvx4));
assign N81wx4 = (~(H3wvx4 & haddr_o[13]));
assign T8jvx4 = (I4zvx4 ? B91wx4 : vis_psp_o[11]);
assign M8jvx4 = (P4zvx4 ? B91wx4 : vis_msp_o[11]);
assign F8jvx4 = (Meyvx4 ? B91wx4 : vis_r14_o[13]);
assign Y7jvx4 = (Teyvx4 ? B91wx4 : vis_r12_o[13]);
assign R7jvx4 = (Afyvx4 ? B91wx4 : vis_r7_o[13]);
assign K7jvx4 = (Hfyvx4 ? B91wx4 : vis_r6_o[13]);
assign D7jvx4 = (Ofyvx4 ? B91wx4 : vis_r5_o[13]);
assign W6jvx4 = (Vfyvx4 ? B91wx4 : vis_r4_o[13]);
assign P6jvx4 = (Feyvx4 ? B91wx4 : vis_r11_o[13]);
assign I6jvx4 = (Ydyvx4 ? B91wx4 : vis_r10_o[13]);
assign B6jvx4 = (Rdyvx4 ? B91wx4 : vis_r9_o[13]);
assign U5jvx4 = (Kdyvx4 ? B91wx4 : vis_r8_o[13]);
assign N5jvx4 = (Ddyvx4 ? B91wx4 : vis_r3_o[13]);
assign G5jvx4 = (Wcyvx4 ? B91wx4 : vis_r2_o[13]);
assign Z4jvx4 = (Siqvx4 ? B91wx4 : vis_r1_o[13]);
assign S4jvx4 = (Xppvx4 ? B91wx4 : vis_r0_o[13]);
assign B91wx4 = (~(I91wx4 & P91wx4));
assign P91wx4 = (W91wx4 & Da1wx4);
assign Da1wx4 = (~(Ka1wx4 & Ra1wx4));
assign Ka1wx4 = (E8bvx4 & X8zvx4);
assign W91wx4 = (~(Bpzvx4 | Ya1wx4));
assign I91wx4 = (Fb1wx4 & Mb1wx4);
assign Fb1wx4 = (Tb1wx4 & Ac1wx4);
assign Ac1wx4 = (~(Dmh2z4[13] & Lhyvx4));
assign Tb1wx4 = (Shyvx4 | Hc1wx4);
assign L4jvx4 = (~(Oc1wx4 & Vc1wx4));
assign Vc1wx4 = (~(Cfdvx4 & F2pvx4));
assign Oc1wx4 = (Cd1wx4 & Jd1wx4);
assign Jd1wx4 = (~(vis_pc_o[11] & W0pvx4));
assign Cd1wx4 = (R1pvx4 | Cqovx4);
assign E4jvx4 = (I4zvx4 ? Qd1wx4 : vis_psp_o[10]);
assign X3jvx4 = (P4zvx4 ? Qd1wx4 : vis_msp_o[10]);
assign Q3jvx4 = (Meyvx4 ? Qd1wx4 : vis_r14_o[12]);
assign J3jvx4 = (Teyvx4 ? Qd1wx4 : vis_r12_o[12]);
assign C3jvx4 = (Afyvx4 ? Qd1wx4 : vis_r7_o[12]);
assign V2jvx4 = (Hfyvx4 ? Qd1wx4 : vis_r6_o[12]);
assign O2jvx4 = (Ofyvx4 ? Qd1wx4 : vis_r5_o[12]);
assign H2jvx4 = (Vfyvx4 ? Qd1wx4 : vis_r4_o[12]);
assign A2jvx4 = (Feyvx4 ? Qd1wx4 : vis_r11_o[12]);
assign T1jvx4 = (Ydyvx4 ? Qd1wx4 : vis_r10_o[12]);
assign M1jvx4 = (Rdyvx4 ? Qd1wx4 : vis_r9_o[12]);
assign F1jvx4 = (Kdyvx4 ? Qd1wx4 : vis_r8_o[12]);
assign Y0jvx4 = (Ddyvx4 ? Qd1wx4 : vis_r3_o[12]);
assign R0jvx4 = (Wcyvx4 ? Qd1wx4 : vis_r2_o[12]);
assign K0jvx4 = (Siqvx4 ? Qd1wx4 : vis_r1_o[12]);
assign D0jvx4 = (Xppvx4 ? Qd1wx4 : vis_r0_o[12]);
assign Qd1wx4 = (~(Xd1wx4 & Ee1wx4));
assign Ee1wx4 = (Le1wx4 & Se1wx4);
assign Se1wx4 = (Shyvx4 | Ze1wx4);
assign Le1wx4 = (Gf1wx4 & Egzvx4);
assign Gf1wx4 = (~(Dmh2z4[12] & Lhyvx4));
assign Xd1wx4 = (Nf1wx4 & Uf1wx4);
assign Nf1wx4 = (T6bvx4 ? Ig1wx4 : Bg1wx4);
assign Ig1wx4 = (Pg1wx4 ? Alzvx4 : Tkzvx4);
assign Bg1wx4 = (Olzvx4 | Pg1wx4);
assign Wzivx4 = (~(Wg1wx4 & Dh1wx4));
assign Dh1wx4 = (~(Rddvx4 & F2pvx4));
assign Wg1wx4 = (Kh1wx4 & Rh1wx4);
assign Rh1wx4 = (R1pvx4 | Owovx4);
assign Owovx4 = (Yh1wx4 & Fi1wx4);
assign Fi1wx4 = (~(Gzvvx4 & Axnvx4));
assign Yh1wx4 = (Mi1wx4 & Ti1wx4);
assign Ti1wx4 = (~(Ykh2z4[10] & Mrsvx4));
assign Mi1wx4 = (~(Dmh2z4[11] & K1wvx4));
assign Kh1wx4 = (~(vis_pc_o[10] & W0pvx4));
assign Pzivx4 = (I4zvx4 ? Aj1wx4 : vis_psp_o[9]);
assign Izivx4 = (P4zvx4 ? Aj1wx4 : vis_msp_o[9]);
assign Bzivx4 = (Meyvx4 ? Aj1wx4 : vis_r14_o[11]);
assign Uyivx4 = (Teyvx4 ? Aj1wx4 : vis_r12_o[11]);
assign Nyivx4 = (Afyvx4 ? Aj1wx4 : vis_r7_o[11]);
assign Gyivx4 = (Hfyvx4 ? Aj1wx4 : vis_r6_o[11]);
assign Zxivx4 = (Ofyvx4 ? Aj1wx4 : vis_r5_o[11]);
assign Sxivx4 = (Vfyvx4 ? Aj1wx4 : vis_r4_o[11]);
assign Lxivx4 = (Feyvx4 ? Aj1wx4 : vis_r11_o[11]);
assign Exivx4 = (Ydyvx4 ? Aj1wx4 : vis_r10_o[11]);
assign Xwivx4 = (Rdyvx4 ? Aj1wx4 : vis_r9_o[11]);
assign Qwivx4 = (Kdyvx4 ? Aj1wx4 : vis_r8_o[11]);
assign Jwivx4 = (Ddyvx4 ? Aj1wx4 : vis_r3_o[11]);
assign Cwivx4 = (Wcyvx4 ? Aj1wx4 : vis_r2_o[11]);
assign Vvivx4 = (Siqvx4 ? Aj1wx4 : vis_r1_o[11]);
assign Ovivx4 = (Xppvx4 ? Aj1wx4 : vis_r0_o[11]);
assign Aj1wx4 = (~(Hj1wx4 & Oj1wx4));
assign Oj1wx4 = (Vj1wx4 & Ck1wx4);
assign Ck1wx4 = (~(Jk1wx4 & Qk1wx4));
assign Jk1wx4 = (I5bvx4 & X8zvx4);
assign Vj1wx4 = (~(Bpzvx4 | Xk1wx4));
assign Hj1wx4 = (El1wx4 & Ll1wx4);
assign El1wx4 = (Sl1wx4 & Zl1wx4);
assign Zl1wx4 = (~(Dmh2z4[11] & Lhyvx4));
assign Sl1wx4 = (Shyvx4 | Gm1wx4);
assign Hvivx4 = (~(Nm1wx4 & Um1wx4));
assign Um1wx4 = (~(Gcdvx4 & F2pvx4));
assign Nm1wx4 = (Bn1wx4 & In1wx4);
assign In1wx4 = (~(vis_pc_o[9] & W0pvx4));
assign Bn1wx4 = (R1pvx4 | Jxovx4);
assign Avivx4 = (I4zvx4 ? Pn1wx4 : vis_psp_o[8]);
assign Tuivx4 = (P4zvx4 ? Pn1wx4 : vis_msp_o[8]);
assign Muivx4 = (Meyvx4 ? Pn1wx4 : vis_r14_o[10]);
assign Fuivx4 = (Teyvx4 ? Pn1wx4 : vis_r12_o[10]);
assign Ytivx4 = (Afyvx4 ? Pn1wx4 : vis_r7_o[10]);
assign Rtivx4 = (Hfyvx4 ? Pn1wx4 : vis_r6_o[10]);
assign Ktivx4 = (Ofyvx4 ? Pn1wx4 : vis_r5_o[10]);
assign Dtivx4 = (Vfyvx4 ? Pn1wx4 : vis_r4_o[10]);
assign Wsivx4 = (Feyvx4 ? Pn1wx4 : vis_r11_o[10]);
assign Psivx4 = (Ydyvx4 ? Pn1wx4 : vis_r10_o[10]);
assign Isivx4 = (Rdyvx4 ? Pn1wx4 : vis_r9_o[10]);
assign Bsivx4 = (Kdyvx4 ? Pn1wx4 : vis_r8_o[10]);
assign Urivx4 = (Ddyvx4 ? Pn1wx4 : vis_r3_o[10]);
assign Nrivx4 = (Wcyvx4 ? Pn1wx4 : vis_r2_o[10]);
assign Grivx4 = (Siqvx4 ? Pn1wx4 : vis_r1_o[10]);
assign Zqivx4 = (Xppvx4 ? Pn1wx4 : vis_r0_o[10]);
assign Pn1wx4 = (~(Wn1wx4 & Do1wx4));
assign Sqivx4 = (Ro1wx4 ? Ko1wx4 : Oy8vx4);
assign Ro1wx4 = (Yo1wx4 & hready_i);
assign Yo1wx4 = (~(Fp1wx4 & Mp1wx4));
assign Mp1wx4 = (~(Tp1wx4 & Aq1wx4));
assign Fp1wx4 = (Hq1wx4 | Jrnvx4);
assign Ko1wx4 = (Mtqvx4 ? Qrnvx4 : Oq1wx4);
assign Oq1wx4 = (!Vq1wx4);
assign Lqivx4 = (I4zvx4 ? Cr1wx4 : vis_psp_o[0]);
assign Eqivx4 = (P4zvx4 ? Cr1wx4 : vis_msp_o[0]);
assign Xpivx4 = (Meyvx4 ? Cr1wx4 : vis_r14_o[2]);
assign Qpivx4 = (Teyvx4 ? Cr1wx4 : vis_r12_o[2]);
assign Jpivx4 = (Afyvx4 ? Cr1wx4 : vis_r7_o[2]);
assign Cpivx4 = (Hfyvx4 ? Cr1wx4 : vis_r6_o[2]);
assign Voivx4 = (Ofyvx4 ? Cr1wx4 : vis_r5_o[2]);
assign Ooivx4 = (Vfyvx4 ? Cr1wx4 : vis_r4_o[2]);
assign Hoivx4 = (Feyvx4 ? Cr1wx4 : vis_r11_o[2]);
assign Aoivx4 = (Ydyvx4 ? Cr1wx4 : vis_r10_o[2]);
assign Tnivx4 = (Rdyvx4 ? Cr1wx4 : vis_r9_o[2]);
assign Mnivx4 = (Kdyvx4 ? Cr1wx4 : vis_r8_o[2]);
assign Fnivx4 = (Ddyvx4 ? Cr1wx4 : vis_r3_o[2]);
assign Ymivx4 = (Wcyvx4 ? Cr1wx4 : vis_r2_o[2]);
assign Rmivx4 = (Siqvx4 ? Cr1wx4 : vis_r1_o[2]);
assign Kmivx4 = (Xppvx4 ? Cr1wx4 : vis_r0_o[2]);
assign Cr1wx4 = (~(Zluvx4 & Jr1wx4));
assign Dmivx4 = (~(Qr1wx4 & Xr1wx4));
assign Xr1wx4 = (Es1wx4 & Ls1wx4);
assign Ls1wx4 = (R1pvx4 | Xxovx4);
assign Xxovx4 = (Ss1wx4 & Zs1wx4);
assign Zs1wx4 = (~(Gzvvx4 & Konvx4));
assign Ss1wx4 = (Gt1wx4 & Nt1wx4);
assign Nt1wx4 = (~(Ykh2z4[8] & Mrsvx4));
assign Gt1wx4 = (~(Dmh2z4[9] & K1wvx4));
assign Es1wx4 = (~(Oy8vx4 & P0pvx4));
assign Qr1wx4 = (Ut1wx4 & Bu1wx4);
assign Bu1wx4 = (~(vis_pc_o[8] & W0pvx4));
assign Ut1wx4 = (~(Wadvx4 & F2pvx4));
assign Wlivx4 = (I4zvx4 ? Iu1wx4 : vis_psp_o[7]);
assign Plivx4 = (P4zvx4 ? Iu1wx4 : vis_msp_o[7]);
assign P4zvx4 = (!Pu1wx4);
assign Ilivx4 = (Meyvx4 ? Iu1wx4 : vis_r14_o[9]);
assign Blivx4 = (Teyvx4 ? Iu1wx4 : vis_r12_o[9]);
assign Teyvx4 = (!Wu1wx4);
assign Ukivx4 = (Afyvx4 ? Iu1wx4 : vis_r7_o[9]);
assign Afyvx4 = (!Dv1wx4);
assign Nkivx4 = (Hfyvx4 ? Iu1wx4 : vis_r6_o[9]);
assign Gkivx4 = (Ofyvx4 ? Iu1wx4 : vis_r5_o[9]);
assign Ofyvx4 = (!Kv1wx4);
assign Zjivx4 = (Vfyvx4 ? Iu1wx4 : vis_r4_o[9]);
assign Vfyvx4 = (!Rv1wx4);
assign Sjivx4 = (Feyvx4 ? Iu1wx4 : vis_r11_o[9]);
assign Feyvx4 = (!Yv1wx4);
assign Ljivx4 = (Ydyvx4 ? Iu1wx4 : vis_r10_o[9]);
assign Ejivx4 = (Rdyvx4 ? Iu1wx4 : vis_r9_o[9]);
assign Rdyvx4 = (!Fw1wx4);
assign Xiivx4 = (Kdyvx4 ? Iu1wx4 : vis_r8_o[9]);
assign Kdyvx4 = (!Mw1wx4);
assign Qiivx4 = (Ddyvx4 ? Iu1wx4 : vis_r3_o[9]);
assign Ddyvx4 = (!Tw1wx4);
assign Jiivx4 = (Wcyvx4 ? Iu1wx4 : vis_r2_o[9]);
assign Ciivx4 = (Siqvx4 ? Iu1wx4 : vis_r1_o[9]);
assign Siqvx4 = (!Ax1wx4);
assign Vhivx4 = (Xppvx4 ? Iu1wx4 : vis_r0_o[9]);
assign Xppvx4 = (!Hx1wx4);
assign Iu1wx4 = (~(Vq1wx4 & Ox1wx4));
assign Ohivx4 = (~(Vx1wx4 & Cy1wx4));
assign Cy1wx4 = (~(M9dvx4 & F2pvx4));
assign Vx1wx4 = (Jy1wx4 & Qy1wx4);
assign Qy1wx4 = (R1pvx4 | Z6ovx4);
assign Z6ovx4 = (Xy1wx4 & Ez1wx4);
assign Ez1wx4 = (~(Gzvvx4 & Ronvx4));
assign Xy1wx4 = (Lz1wx4 & Sz1wx4);
assign Sz1wx4 = (~(Ykh2z4[7] & Mrsvx4));
assign Lz1wx4 = (~(Dmh2z4[8] & K1wvx4));
assign Jy1wx4 = (~(vis_pc_o[7] & W0pvx4));
assign Hhivx4 = (I4zvx4 ? Zz1wx4 : vis_psp_o[6]);
assign I4zvx4 = (!G02wx4);
assign Ahivx4 = (Pu1wx4 ? vis_msp_o[6] : Zz1wx4);
assign Tgivx4 = (Meyvx4 ? Zz1wx4 : vis_r14_o[8]);
assign Mgivx4 = (Wu1wx4 ? vis_r12_o[8] : Zz1wx4);
assign Fgivx4 = (Dv1wx4 ? vis_r7_o[8] : Zz1wx4);
assign Yfivx4 = (Hfyvx4 ? Zz1wx4 : vis_r6_o[8]);
assign Rfivx4 = (Kv1wx4 ? vis_r5_o[8] : Zz1wx4);
assign Kfivx4 = (Rv1wx4 ? vis_r4_o[8] : Zz1wx4);
assign Dfivx4 = (Yv1wx4 ? vis_r11_o[8] : Zz1wx4);
assign Weivx4 = (Ydyvx4 ? Zz1wx4 : vis_r10_o[8]);
assign Peivx4 = (Fw1wx4 ? vis_r9_o[8] : Zz1wx4);
assign Ieivx4 = (Mw1wx4 ? vis_r8_o[8] : Zz1wx4);
assign Beivx4 = (Tw1wx4 ? vis_r3_o[8] : Zz1wx4);
assign Udivx4 = (Wcyvx4 ? Zz1wx4 : vis_r2_o[8]);
assign Ndivx4 = (Ax1wx4 ? vis_r1_o[8] : Zz1wx4);
assign Gdivx4 = (Hx1wx4 ? vis_r0_o[8] : Zz1wx4);
assign Zz1wx4 = (~(N02wx4 & U02wx4));
assign U02wx4 = (B12wx4 & I12wx4);
assign I12wx4 = (Shyvx4 | P12wx4);
assign B12wx4 = (W12wx4 & Egzvx4);
assign W12wx4 = (~(Dmh2z4[8] & Lhyvx4));
assign N02wx4 = (D22wx4 & K22wx4);
assign D22wx4 = (Y3bvx4 ? Y22wx4 : R22wx4);
assign Y22wx4 = (F32wx4 ? Alzvx4 : Tkzvx4);
assign R22wx4 = (Olzvx4 | F32wx4);
assign Zcivx4 = (~(M32wx4 & T32wx4));
assign T32wx4 = (~(Jjdvx4 & F2pvx4));
assign M32wx4 = (A42wx4 & H42wx4);
assign H42wx4 = (~(H3wvx4 & haddr_o[15]));
assign haddr_o[15] = (~(O42wx4 & V42wx4));
assign V42wx4 = (~(Gzvvx4 & Yvnvx4));
assign O42wx4 = (C52wx4 & J52wx4);
assign J52wx4 = (~(Ykh2z4[14] & Mrsvx4));
assign C52wx4 = (~(Dmh2z4[15] & K1wvx4));
assign A42wx4 = (~(vis_pc_o[14] & W0pvx4));
assign Scivx4 = (G02wx4 ? vis_psp_o[13] : Q52wx4);
assign Lcivx4 = (Pu1wx4 ? vis_msp_o[13] : Q52wx4);
assign Ecivx4 = (Meyvx4 ? Q52wx4 : vis_r14_o[15]);
assign Xbivx4 = (Wu1wx4 ? vis_r12_o[15] : Q52wx4);
assign Qbivx4 = (Dv1wx4 ? vis_r7_o[15] : Q52wx4);
assign Jbivx4 = (Hfyvx4 ? Q52wx4 : vis_r6_o[15]);
assign Cbivx4 = (Kv1wx4 ? vis_r5_o[15] : Q52wx4);
assign Vaivx4 = (Rv1wx4 ? vis_r4_o[15] : Q52wx4);
assign Oaivx4 = (Yv1wx4 ? vis_r11_o[15] : Q52wx4);
assign Haivx4 = (Ydyvx4 ? Q52wx4 : vis_r10_o[15]);
assign Aaivx4 = (Fw1wx4 ? vis_r9_o[15] : Q52wx4);
assign T9ivx4 = (Mw1wx4 ? vis_r8_o[15] : Q52wx4);
assign M9ivx4 = (Tw1wx4 ? vis_r3_o[15] : Q52wx4);
assign F9ivx4 = (Wcyvx4 ? Q52wx4 : vis_r2_o[15]);
assign Y8ivx4 = (Ax1wx4 ? vis_r1_o[15] : Q52wx4);
assign R8ivx4 = (Hx1wx4 ? vis_r0_o[15] : Q52wx4);
assign Q52wx4 = (~(X52wx4 & E62wx4));
assign E62wx4 = (L62wx4 & S62wx4);
assign S62wx4 = (Shyvx4 | Z62wx4);
assign L62wx4 = (G72wx4 & Egzvx4);
assign G72wx4 = (~(Dmh2z4[15] & Lhyvx4));
assign X52wx4 = (N72wx4 & U72wx4);
assign N72wx4 = (Abbvx4 ? I82wx4 : B82wx4);
assign I82wx4 = (P82wx4 ? Alzvx4 : Tkzvx4);
assign B82wx4 = (Olzvx4 | P82wx4);
assign K8ivx4 = (~(W82wx4 & D92wx4));
assign D92wx4 = (~(Tudvx4 & F2pvx4));
assign W82wx4 = (K92wx4 & R92wx4);
assign R92wx4 = (~(vis_pc_o[22] & W0pvx4));
assign K92wx4 = (R1pvx4 | Y92wx4);
assign D8ivx4 = (G02wx4 ? vis_psp_o[21] : Fa2wx4);
assign G02wx4 = (Ma2wx4 | Ta2wx4);
assign W7ivx4 = (Pu1wx4 ? vis_msp_o[21] : Fa2wx4);
assign Pu1wx4 = (Ma2wx4 | O7evx4);
assign Ma2wx4 = (~(Ab2wx4 & Hb2wx4));
assign Ab2wx4 = (~(Ob2wx4 | Vb2wx4));
assign P7ivx4 = (Meyvx4 ? Fa2wx4 : vis_r14_o[23]);
assign Meyvx4 = (Cc2wx4 & Jc2wx4);
assign I7ivx4 = (Wu1wx4 ? vis_r12_o[23] : Fa2wx4);
assign Wu1wx4 = (~(Qc2wx4 & Cc2wx4));
assign Qc2wx4 = (Xc2wx4 & Ed2wx4);
assign B7ivx4 = (Dv1wx4 ? vis_r7_o[23] : Fa2wx4);
assign Dv1wx4 = (~(Ld2wx4 & Sd2wx4));
assign Ld2wx4 = (Zd2wx4 & Ge2wx4);
assign U6ivx4 = (Hfyvx4 ? Fa2wx4 : vis_r6_o[23]);
assign Hfyvx4 = (Cc2wx4 & Sd2wx4);
assign N6ivx4 = (Kv1wx4 ? vis_r5_o[23] : Fa2wx4);
assign Kv1wx4 = (~(Ne2wx4 & Hb2wx4));
assign Ne2wx4 = (~(Ed2wx4 | Vb2wx4));
assign G6ivx4 = (Rv1wx4 ? vis_r4_o[23] : Fa2wx4);
assign Rv1wx4 = (~(Ue2wx4 & Cc2wx4));
assign Cc2wx4 = (~(Ge2wx4 | Vb2wx4));
assign Ue2wx4 = (Xc2wx4 & Ob2wx4);
assign Z5ivx4 = (Yv1wx4 ? vis_r11_o[23] : Fa2wx4);
assign Yv1wx4 = (~(Bf2wx4 & Jc2wx4));
assign S5ivx4 = (Ydyvx4 ? Fa2wx4 : vis_r10_o[23]);
assign Ydyvx4 = (Jc2wx4 & If2wx4);
assign Jc2wx4 = (~(Ob2wx4 | Xc2wx4));
assign L5ivx4 = (Fw1wx4 ? vis_r9_o[23] : Fa2wx4);
assign Fw1wx4 = (~(Pf2wx4 & Hb2wx4));
assign Pf2wx4 = (~(Zd2wx4 | Ob2wx4));
assign E5ivx4 = (Mw1wx4 ? vis_r8_o[23] : Fa2wx4);
assign Mw1wx4 = (~(Wf2wx4 & Xc2wx4));
assign Wf2wx4 = (If2wx4 & Ed2wx4);
assign X4ivx4 = (Tw1wx4 ? vis_r3_o[23] : Fa2wx4);
assign Tw1wx4 = (~(Bf2wx4 & Sd2wx4));
assign Bf2wx4 = (Vb2wx4 & Ge2wx4);
assign Q4ivx4 = (Wcyvx4 ? Fa2wx4 : vis_r2_o[23]);
assign Wcyvx4 = (Sd2wx4 & If2wx4);
assign Sd2wx4 = (~(Ed2wx4 | Xc2wx4));
assign J4ivx4 = (Ax1wx4 ? vis_r1_o[23] : Fa2wx4);
assign Ax1wx4 = (~(Dg2wx4 & Hb2wx4));
assign Hb2wx4 = (Xc2wx4 & Ge2wx4);
assign Dg2wx4 = (~(Ed2wx4 | Zd2wx4));
assign Ed2wx4 = (!Ob2wx4);
assign C4ivx4 = (Hx1wx4 ? vis_r0_o[23] : Fa2wx4);
assign Hx1wx4 = (~(Kg2wx4 & Xc2wx4));
assign Xc2wx4 = (Rg2wx4 & Yg2wx4);
assign Rg2wx4 = (Fh2wx4 & hready_i);
assign Kg2wx4 = (Ob2wx4 & If2wx4);
assign If2wx4 = (~(Ge2wx4 | Zd2wx4));
assign Zd2wx4 = (!Vb2wx4);
assign Vb2wx4 = (Mh2wx4 & Th2wx4);
assign Th2wx4 = (Ai2wx4 & Hi2wx4);
assign Hi2wx4 = (~(Wv9vx4 & Oi2wx4));
assign Ai2wx4 = (~(Nt8vx4 & Vi2wx4));
assign Mh2wx4 = (Cj2wx4 & Jj2wx4);
assign Jj2wx4 = (~(Tjh2z4[2] & Qj2wx4));
assign Ge2wx4 = (~(Xj2wx4 & Ek2wx4));
assign Ek2wx4 = (Lk2wx4 & Sk2wx4);
assign Sk2wx4 = (~(Tjh2z4[0] & Qj2wx4));
assign Lk2wx4 = (~(Ot9vx4 & Oi2wx4));
assign Xj2wx4 = (Zk2wx4 & Gl2wx4);
assign Gl2wx4 = (~(Xq8vx4 & Vi2wx4));
assign Ob2wx4 = (Nl2wx4 & Ul2wx4);
assign Ul2wx4 = (Bm2wx4 & Im2wx4);
assign Im2wx4 = (~(Bx9vx4 & Oi2wx4));
assign Bm2wx4 = (~(Vu8vx4 & Vi2wx4));
assign Nl2wx4 = (Cj2wx4 & Pm2wx4);
assign Pm2wx4 = (~(Tjh2z4[3] & Qj2wx4));
assign Cj2wx4 = (Wm2wx4 & Zk2wx4);
assign Zk2wx4 = (Dn2wx4 & Fh2wx4);
assign Fh2wx4 = (~(Kn2wx4 & Rn2wx4));
assign Rn2wx4 = (Yn2wx4 & Fo2wx4);
assign Fo2wx4 = (Mo2wx4 & To2wx4);
assign To2wx4 = (~(Ap2wx4 & Huqvx4));
assign Ap2wx4 = (~(Hp2wx4 | Nggvx4));
assign Mo2wx4 = (Op2wx4 & Vp2wx4);
assign Yn2wx4 = (Cq2wx4 & Jq2wx4);
assign Jq2wx4 = (~(U9gvx4 & Qq2wx4));
assign Qq2wx4 = (~(Xq2wx4 & Er2wx4));
assign Er2wx4 = (Lr2wx4 | Sr2wx4);
assign Xq2wx4 = (~(Zr2wx4 | Gs2wx4));
assign Zr2wx4 = (Ns2wx4 & Kzxvx4);
assign Ns2wx4 = (~(Us2wx4 | Mj8vx4));
assign Cq2wx4 = (Bt2wx4 & It2wx4);
assign It2wx4 = (~(Pt2wx4 & Eiqvx4));
assign Pt2wx4 = (~(Wt2wx4 | Vdgvx4));
assign Bt2wx4 = (~(Du2wx4 & R7qvx4));
assign Du2wx4 = (~(Ku2wx4 & Ru2wx4));
assign Ru2wx4 = (~(Yu2wx4 & Fv2wx4));
assign Yu2wx4 = (~(Mv2wx4 | Tv2wx4));
assign Ku2wx4 = (~(Aw2wx4 & O9qvx4));
assign Aw2wx4 = (Vdgvx4 & Hw2wx4);
assign Kn2wx4 = (Ow2wx4 & Vw2wx4);
assign Vw2wx4 = (Cx2wx4 & Jx2wx4);
assign Jx2wx4 = (~(Qx2wx4 & Xx2wx4));
assign Cx2wx4 = (Ey2wx4 & Ly2wx4);
assign Ly2wx4 = (~(Sy2wx4 & Zy2wx4));
assign Zy2wx4 = (~(Gz2wx4 & Nz2wx4));
assign Nz2wx4 = (~(Uz2wx4 & Zrvvx4));
assign Uz2wx4 = (~(B03wx4 & I03wx4));
assign I03wx4 = (~(P03wx4 & R7qvx4));
assign Gz2wx4 = (~(W03wx4 | D13wx4));
assign W03wx4 = (K13wx4 & Ucqvx4);
assign K13wx4 = (R13wx4 & Mcgvx4);
assign Ey2wx4 = (~(Y13wx4 & F23wx4));
assign F23wx4 = (~(M23wx4 & T23wx4));
assign T23wx4 = (A33wx4 & H33wx4);
assign A33wx4 = (O33wx4 | S4xvx4);
assign M23wx4 = (~(V33wx4 | C43wx4));
assign C43wx4 = (~(J43wx4 | U0ovx4));
assign V33wx4 = (B1ovx4 ? X43wx4 : Q43wx4);
assign Ow2wx4 = (E53wx4 & L53wx4);
assign L53wx4 = (F3ovx4 ? Z53wx4 : S53wx4);
assign Z53wx4 = (G63wx4 & N63wx4);
assign N63wx4 = (~(U63wx4 & B73wx4));
assign G63wx4 = (I73wx4 & P73wx4);
assign P73wx4 = (~(W73wx4 & D83wx4));
assign W73wx4 = (Wkxvx4 & Zrvvx4);
assign I73wx4 = (~(K83wx4 & Xx2wx4));
assign K83wx4 = (Hw2wx4 & S4xvx4);
assign S53wx4 = (R83wx4 & Y83wx4);
assign Y83wx4 = (~(F93wx4 & D83wx4));
assign F93wx4 = (~(M93wx4 | T93wx4));
assign R83wx4 = (~(Wdxvx4 & Huqvx4));
assign E53wx4 = (Aa3wx4 & Ha3wx4);
assign Ha3wx4 = (~(T1xvx4 & Eznvx4));
assign Aa3wx4 = (~(P5yvx4 & Wdxvx4));
assign Dn2wx4 = (~(Ccovx4 | A0zvx4));
assign Fa2wx4 = (~(Oa3wx4 & Va3wx4));
assign V3ivx4 = (Z9zvx4 ? vis_apsr_o[3] : Cb3wx4);
assign Z9zvx4 = (~(Jb3wx4 & hready_i));
assign Jb3wx4 = (~(Qb3wx4 & Wspvx4));
assign Cb3wx4 = (~(Xb3wx4 & Ec3wx4));
assign Ec3wx4 = (~(H3pvx4 & Lc3wx4));
assign Lc3wx4 = (!R5zvx4);
assign H3pvx4 = (!X4pvx4);
assign Xb3wx4 = (Sc3wx4 & Zc3wx4);
assign Zc3wx4 = (Grpvx4 | Gd3wx4);
assign Grpvx4 = (!Wspvx4);
assign Wspvx4 = (X4pvx4 & Ktpvx4);
assign X4pvx4 = (Hq1wx4 | Mtqvx4);
assign Sc3wx4 = (Ktpvx4 | Nd3wx4);
assign Ktpvx4 = (!K0qvx4);
assign K0qvx4 = (Ud3wx4 & Kryvx4);
assign O3ivx4 = (~(Be3wx4 & Ie3wx4));
assign Ie3wx4 = (Pe3wx4 & We3wx4);
assign We3wx4 = (~(vis_apsr_o[3] & P0pvx4));
assign P0pvx4 = (~(F2pvx4 | Vp2wx4));
assign Pe3wx4 = (~(W0pvx4 & vis_pc_o[30]));
assign W0pvx4 = (Df3wx4 & P6xvx4);
assign Be3wx4 = (Kf3wx4 & Rf3wx4);
assign Rf3wx4 = (~(H3wvx4 & haddr_o[31]));
assign H3wvx4 = (!R1pvx4);
assign R1pvx4 = (~(Df3wx4 & Yf3wx4));
assign Yf3wx4 = (~(Fg3wx4 & Mg3wx4));
assign Mg3wx4 = (Gjxvx4 | Dbgvx4);
assign Fg3wx4 = (Tg3wx4 & Jhxvx4);
assign Tg3wx4 = (~(Ah3wx4 & Zrvvx4));
assign Ah3wx4 = (~(Hh3wx4 & Lcpvx4));
assign Kf3wx4 = (~(D6evx4 & F2pvx4));
assign F2pvx4 = (!Df3wx4);
assign Df3wx4 = (hready_i & Oh3wx4);
assign Oh3wx4 = (~(Vh3wx4 & Ci3wx4));
assign Ci3wx4 = (Ji3wx4 & Qi3wx4);
assign Qi3wx4 = (Xi3wx4 & Ej3wx4);
assign Xi3wx4 = (~(Lj3wx4 & Sj3wx4));
assign Sj3wx4 = (~(Zj3wx4 | F3ovx4));
assign Lj3wx4 = (Liqvx4 & P03wx4);
assign Ji3wx4 = (Gk3wx4 & Nk3wx4);
assign Nk3wx4 = (~(Uk3wx4 & Lxwvx4));
assign Uk3wx4 = (Ukpvx4 & Cf9vx4);
assign Gk3wx4 = (~(B4zvx4 & Bl3wx4));
assign Vh3wx4 = (Il3wx4 & Pl3wx4);
assign Pl3wx4 = (Wl3wx4 & Dm3wx4);
assign Dm3wx4 = (~(Km3wx4 & O4ovx4));
assign Km3wx4 = (~(Rm3wx4 & Ym3wx4));
assign Ym3wx4 = (Fn3wx4 & Mn3wx4);
assign Fn3wx4 = (~(Tn3wx4 & Sjwvx4));
assign Tn3wx4 = (V1yvx4 & Ao3wx4);
assign Ao3wx4 = (~(Hh3wx4 & Ho3wx4));
assign Rm3wx4 = (Oo3wx4 & Vo3wx4);
assign Vo3wx4 = (~(Cp3wx4 & Kg9vx4));
assign Oo3wx4 = (~(Jp3wx4 & Qp3wx4));
assign Wl3wx4 = (Xp3wx4 | Jppvx4);
assign Il3wx4 = (~(Eq3wx4 | Lq3wx4));
assign Lq3wx4 = (!Nbyvx4);
assign Eq3wx4 = (M3ovx4 ? Ohpvx4 : Sq3wx4);
assign Ohpvx4 = (!Zq3wx4);
assign Sq3wx4 = (T1xvx4 & Us2wx4);
assign H3ivx4 = (Ih8vx4 ? Nr3wx4 : Gr3wx4);
assign Nr3wx4 = (~(Ur3wx4 & Bs3wx4));
assign Bs3wx4 = (Is3wx4 & Mcgvx4);
assign Is3wx4 = (Xx2wx4 & Ps3wx4);
assign Ur3wx4 = (Ws3wx4 & Ffqvx4);
assign Gr3wx4 = (~(Dt3wx4 & Kt3wx4));
assign Kt3wx4 = (Rt3wx4 & Maovx4);
assign Maovx4 = (!L7uvx4);
assign L7uvx4 = (~(Yt3wx4 | K7xvx4));
assign Rt3wx4 = (~(rxev_i | txev_o));
assign txev_o = (~(Fu3wx4 | Mu3wx4));
assign Fu3wx4 = (~(Vdgvx4 & Ps3wx4));
assign Dt3wx4 = (Tu3wx4 & Vbovx4);
assign Tu3wx4 = (~(Vogvx4 & Av3wx4));
assign Av3wx4 = (~(Hv3wx4 & Ov3wx4));
assign Ov3wx4 = (Vv3wx4 & Cw3wx4);
assign Cw3wx4 = (Jw3wx4 & Qw3wx4);
assign Qw3wx4 = (Xw3wx4 & Ex3wx4);
assign Ex3wx4 = (~(Lx3wx4 & Pmvvx4));
assign Lx3wx4 = (~(Sx3wx4 | Qsgvx4));
assign Xw3wx4 = (Zx3wx4 & Gy3wx4);
assign Gy3wx4 = (~(D9ovx4 & Ny3wx4));
assign Ny3wx4 = (~(Uy3wx4 & Bz3wx4));
assign Bz3wx4 = (Iz3wx4 & Pz3wx4);
assign Pz3wx4 = (Wz3wx4 & D04wx4);
assign Wz3wx4 = (~(hwdata_o[27] | hwdata_o[28]));
assign Iz3wx4 = (K04wx4 & R04wx4);
assign R04wx4 = (~(hwdata_o[25] | hwdata_o[26]));
assign K04wx4 = (~(Cztvx4 | hwdata_o[24]));
assign Uy3wx4 = (Y04wx4 & F14wx4);
assign F14wx4 = (M14wx4 & T14wx4);
assign T14wx4 = (~(hwdata_o[17] | V4ovx4));
assign M14wx4 = (~(hwdata_o[20] | hwdata_o[18]));
assign Y04wx4 = (A24wx4 & H24wx4);
assign H24wx4 = (~(hwdata_o[16] | hwdata_o[21]));
assign hwdata_o[16] = (!O24wx4);
assign A24wx4 = (~(hwdata_o[22] | hwdata_o[19]));
assign Zx3wx4 = (~(V24wx4 & C34wx4));
assign V24wx4 = (~(Cjvvx4 | Wtgvx4));
assign Cjvvx4 = (J34wx4 & Q34wx4);
assign Q34wx4 = (~(X34wx4 & E44wx4));
assign X34wx4 = (~(Jhxvx4 | J43wx4));
assign Jw3wx4 = (L44wx4 & S44wx4);
assign S44wx4 = (Z44wx4 | T1i2z4[15]);
assign Z44wx4 = (!Syhvx4);
assign L44wx4 = (G54wx4 & N54wx4);
assign N54wx4 = (Ynvvx4 | R3hvx4);
assign Ynvvx4 = (U54wx4 & B64wx4);
assign B64wx4 = (~(I64wx4 & H5uvx4));
assign H5uvx4 = (Irh2z4[0] & F2hvx4);
assign I64wx4 = (Oytvx4 & S0hvx4);
assign Oytvx4 = (P64wx4 & W64wx4);
assign W64wx4 = (D74wx4 & K74wx4);
assign K74wx4 = (R74wx4 & Y74wx4);
assign Y74wx4 = (~(F84wx4 | Irh2z4[7]));
assign F84wx4 = (Irh2z4[8] | Irh2z4[9]);
assign R74wx4 = (~(M84wx4 | Irh2z4[4]));
assign M84wx4 = (Irh2z4[5] | Irh2z4[6]);
assign D74wx4 = (T84wx4 & A94wx4);
assign A94wx4 = (~(H94wx4 | Irh2z4[23]));
assign H94wx4 = (Irh2z4[2] | Irh2z4[3]);
assign T84wx4 = (~(O94wx4 | Irh2z4[20]));
assign O94wx4 = (Irh2z4[21] | Irh2z4[22]);
assign P64wx4 = (V94wx4 & Ca4wx4);
assign Ca4wx4 = (Ja4wx4 & Qa4wx4);
assign Qa4wx4 = (~(Xa4wx4 | Irh2z4[18]));
assign Xa4wx4 = (Irh2z4[19] | Irh2z4[1]);
assign Ja4wx4 = (~(Eb4wx4 | Irh2z4[15]));
assign Eb4wx4 = (Irh2z4[16] | Irh2z4[17]);
assign V94wx4 = (Lb4wx4 & Sb4wx4);
assign Sb4wx4 = (~(Zb4wx4 | Irh2z4[12]));
assign Zb4wx4 = (Irh2z4[13] | Irh2z4[14]);
assign Lb4wx4 = (~(Irh2z4[10] | Irh2z4[11]));
assign U54wx4 = (~(Pmvvx4 & hwdata_o[26]));
assign Pmvvx4 = (Gc4wx4 & Mf8vx4);
assign G54wx4 = (Q5vvx4 | Krgvx4);
assign Q5vvx4 = (Nc4wx4 & Uc4wx4);
assign Uc4wx4 = (J34wx4 | C34wx4);
assign J34wx4 = (~(Bd4wx4 & Id4wx4));
assign Id4wx4 = (~(Mj8vx4 | Vdgvx4));
assign Bd4wx4 = (~(Mu3wx4 | Zj3wx4));
assign Nc4wx4 = (Pd4wx4 & Wd4wx4);
assign Wd4wx4 = (~(De4wx4 & Ke4wx4));
assign Ke4wx4 = (Re4wx4 & C5vvx4);
assign Re4wx4 = (~(Mtqvx4 & Ye4wx4));
assign Mtqvx4 = (Ff4wx4 & Mf4wx4);
assign Mf4wx4 = (Tf4wx4 & Ag4wx4);
assign Ag4wx4 = (~(Mj8vx4 & Hg4wx4));
assign Tf4wx4 = (Vp2wx4 & Og4wx4);
assign Ff4wx4 = (Vg4wx4 & Ch4wx4);
assign Ch4wx4 = (~(Tp1wx4 & Jh4wx4));
assign Jh4wx4 = (~(F3ovx4 | Nggvx4));
assign Tp1wx4 = (P03wx4 & Sy2wx4);
assign De4wx4 = (~(R7qvx4 | Zrvvx4));
assign Pd4wx4 = (~(Qh4wx4 & O4vvx4));
assign Qh4wx4 = (~(Xh4wx4 & Ei4wx4));
assign Ei4wx4 = (Li4wx4 & Si4wx4);
assign Si4wx4 = (~(Zi4wx4 & Gj4wx4));
assign Gj4wx4 = (O9qvx4 & Pcyvx4);
assign Zi4wx4 = (Nj4wx4 & Eznvx4);
assign Li4wx4 = (~(Uj4wx4 & Bk4wx4));
assign Xh4wx4 = (Ik4wx4 & Pk4wx4);
assign Pk4wx4 = (~(Wk4wx4 & Dmgvx4));
assign Wk4wx4 = (~(Zrvvx4 | C5vvx4));
assign Vv3wx4 = (Dl4wx4 & Kl4wx4);
assign Kl4wx4 = (Rl4wx4 & Yl4wx4);
assign Yl4wx4 = (Fm4wx4 | T1i2z4[12]);
assign Fm4wx4 = (!Nzhvx4);
assign Rl4wx4 = (Mm4wx4 & Tm4wx4);
assign Tm4wx4 = (An4wx4 | T1i2z4[14]);
assign An4wx4 = (!Zyhvx4);
assign Mm4wx4 = (Hn4wx4 | T1i2z4[13]);
assign Hn4wx4 = (!Gzhvx4);
assign Dl4wx4 = (On4wx4 & Vn4wx4);
assign Vn4wx4 = (Co4wx4 | T1i2z4[11]);
assign Co4wx4 = (!Uzhvx4);
assign On4wx4 = (Jo4wx4 | T1i2z4[10]);
assign Jo4wx4 = (!B0ivx4);
assign Hv3wx4 = (Qo4wx4 & Xo4wx4);
assign Xo4wx4 = (Ep4wx4 & Lp4wx4);
assign Lp4wx4 = (Sp4wx4 & Zp4wx4);
assign Zp4wx4 = (Gq4wx4 | T1i2z4[7]);
assign Gq4wx4 = (!W0ivx4);
assign Sp4wx4 = (Nq4wx4 & Uq4wx4);
assign Uq4wx4 = (Br4wx4 | T1i2z4[9]);
assign Br4wx4 = (!I0ivx4);
assign Nq4wx4 = (Ir4wx4 | T1i2z4[8]);
assign Ir4wx4 = (!P0ivx4);
assign Ep4wx4 = (Pr4wx4 & Wr4wx4);
assign Wr4wx4 = (Ds4wx4 | T1i2z4[4]);
assign Ds4wx4 = (!R1ivx4);
assign Pr4wx4 = (Ks4wx4 & Rs4wx4);
assign Rs4wx4 = (Ys4wx4 | T1i2z4[6]);
assign Ys4wx4 = (!D1ivx4);
assign Ks4wx4 = (Ft4wx4 | T1i2z4[5]);
assign Ft4wx4 = (!K1ivx4);
assign Qo4wx4 = (Mt4wx4 & Tt4wx4);
assign Tt4wx4 = (Au4wx4 & Hu4wx4);
assign Hu4wx4 = (Ou4wx4 | T1i2z4[1]);
assign Ou4wx4 = (!M2ivx4);
assign Au4wx4 = (Vu4wx4 & Cv4wx4);
assign Cv4wx4 = (Jv4wx4 | T1i2z4[3]);
assign Jv4wx4 = (!Y1ivx4);
assign Vu4wx4 = (Qv4wx4 | T1i2z4[2]);
assign Qv4wx4 = (!F2ivx4);
assign Mt4wx4 = (Xv4wx4 & Ew4wx4);
assign Ew4wx4 = (Lw4wx4 | T1i2z4[0]);
assign Lw4wx4 = (!T2ivx4);
assign Xv4wx4 = (~(Owgvx4 & Sw4wx4));
assign Owgvx4 = (R2vvx4 & Zw4wx4);
assign Zw4wx4 = (~(Gx4wx4 & Nx4wx4));
assign Nx4wx4 = (~(nmi_i & K2vvx4));
assign K2vvx4 = (!Aygvx4);
assign Gx4wx4 = (D2vvx4 & Sw4wx4);
assign D2vvx4 = (~(Cztvx4 & Gc4wx4));
assign Cztvx4 = (!Ux4wx4);
assign R2vvx4 = (~(F3vvx4 & Fsyvx4));
assign Fsyvx4 = (!Vbovx4);
assign A3ivx4 = (!By4wx4);
assign T2ivx4 = (I8ovx4 & Iy4wx4);
assign Iy4wx4 = (~(Py4wx4 & Wy4wx4));
assign Wy4wx4 = (~(irq_i[0] & B8ovx4));
assign B8ovx4 = (!D3i2z4[0]);
assign Py4wx4 = (Dz4wx4 & Kz4wx4);
assign Kz4wx4 = (~(T1i2z4[0] & Rz4wx4));
assign Rz4wx4 = (~(Yz4wx4 & hwdata_o[0]));
assign Dz4wx4 = (~(D9ovx4 & hwdata_o[0]));
assign I8ovx4 = (Taovx4 | Vbovx4);
assign M2ivx4 = (Itvvx4 & F05wx4);
assign F05wx4 = (~(M05wx4 & T05wx4));
assign T05wx4 = (~(irq_i[1] & Btvvx4));
assign Btvvx4 = (!D3i2z4[1]);
assign M05wx4 = (Kuvvx4 & A15wx4);
assign A15wx4 = (~(T1i2z4[1] & H15wx4));
assign H15wx4 = (~(Yz4wx4 & hwdata_o[1]));
assign hwdata_o[1] = (!O15wx4);
assign Kuvvx4 = (V15wx4 | O15wx4);
assign O15wx4 = (~(Pp8vx4 & Htyvx4));
assign Itvvx4 = (Ruvvx4 | Vbovx4);
assign F2ivx4 = (Tiuvx4 & C25wx4);
assign C25wx4 = (~(J25wx4 & Q25wx4));
assign Q25wx4 = (~(irq_i[2] & Miuvx4));
assign Miuvx4 = (!D3i2z4[2]);
assign J25wx4 = (Vjuvx4 & X25wx4);
assign X25wx4 = (~(T1i2z4[2] & E35wx4));
assign E35wx4 = (~(Yz4wx4 & hwdata_o[2]));
assign Vjuvx4 = (V15wx4 | L35wx4);
assign Tiuvx4 = (Ckuvx4 | Vbovx4);
assign Y1ivx4 = (Ufuvx4 & S35wx4);
assign S35wx4 = (~(Z35wx4 & G45wx4));
assign G45wx4 = (~(irq_i[3] & Nfuvx4));
assign Nfuvx4 = (!D3i2z4[3]);
assign Z35wx4 = (N45wx4 & U45wx4);
assign U45wx4 = (~(T1i2z4[3] & B55wx4));
assign B55wx4 = (~(Yz4wx4 & hwdata_o[3]));
assign N45wx4 = (~(D9ovx4 & hwdata_o[3]));
assign Ufuvx4 = (Khuvx4 | Vbovx4);
assign R1ivx4 = (Twuvx4 & I55wx4);
assign I55wx4 = (~(P55wx4 & W55wx4));
assign W55wx4 = (~(irq_i[4] & Mwuvx4));
assign Mwuvx4 = (!D3i2z4[4]);
assign P55wx4 = (D65wx4 & K65wx4);
assign K65wx4 = (~(T1i2z4[4] & R65wx4));
assign R65wx4 = (~(Yz4wx4 & hwdata_o[4]));
assign D65wx4 = (V15wx4 | Jyuvx4);
assign Twuvx4 = (Qyuvx4 | Vbovx4);
assign K1ivx4 = (Ntuvx4 & Y65wx4);
assign Y65wx4 = (~(F75wx4 & M75wx4));
assign M75wx4 = (~(irq_i[5] & Gtuvx4));
assign Gtuvx4 = (!D3i2z4[5]);
assign F75wx4 = (T75wx4 & A85wx4);
assign A85wx4 = (~(T1i2z4[5] & H85wx4));
assign H85wx4 = (~(Yz4wx4 & hwdata_o[5]));
assign T75wx4 = (V15wx4 | Dvuvx4);
assign Ntuvx4 = (Kvuvx4 | Vbovx4);
assign D1ivx4 = (Oquvx4 & O85wx4);
assign O85wx4 = (~(V85wx4 & C95wx4));
assign C95wx4 = (~(irq_i[6] & Hquvx4));
assign Hquvx4 = (!D3i2z4[6]);
assign V85wx4 = (J95wx4 & Q95wx4);
assign Q95wx4 = (~(T1i2z4[6] & X95wx4));
assign X95wx4 = (~(Yz4wx4 & hwdata_o[6]));
assign J95wx4 = (~(D9ovx4 & hwdata_o[6]));
assign Oquvx4 = (Esuvx4 | Vbovx4);
assign W0ivx4 = (Inuvx4 & Ea5wx4);
assign Ea5wx4 = (~(La5wx4 & Sa5wx4));
assign Sa5wx4 = (~(irq_i[7] & Bnuvx4));
assign Bnuvx4 = (!D3i2z4[7]);
assign La5wx4 = (Za5wx4 & Gb5wx4);
assign Gb5wx4 = (~(T1i2z4[7] & Nb5wx4));
assign Nb5wx4 = (~(Yz4wx4 & hwdata_o[7]));
assign Za5wx4 = (V15wx4 | Youvx4);
assign Inuvx4 = (Fpuvx4 | Vbovx4);
assign P0ivx4 = (Dgvvx4 & Ub5wx4);
assign Ub5wx4 = (~(Bc5wx4 & Ic5wx4));
assign Ic5wx4 = (~(irq_i[8] & Wfvvx4));
assign Wfvvx4 = (!D3i2z4[8]);
assign Bc5wx4 = (Fhvvx4 & Pc5wx4);
assign Pc5wx4 = (~(T1i2z4[8] & Wc5wx4));
assign Wc5wx4 = (~(Yz4wx4 & hwdata_o[8]));
assign Fhvvx4 = (V15wx4 | Dd5wx4);
assign Dd5wx4 = (!hwdata_o[8]);
assign hwdata_o[8] = (Yd5wx4 ? Rd5wx4 : Kd5wx4);
assign Dgvvx4 = (Mhvvx4 | Vbovx4);
assign I0ivx4 = (Ldvvx4 & Fe5wx4);
assign Fe5wx4 = (~(Me5wx4 & Te5wx4));
assign Te5wx4 = (~(irq_i[9] & Edvvx4));
assign Edvvx4 = (!D3i2z4[9]);
assign Me5wx4 = (Nevvx4 & Af5wx4);
assign Af5wx4 = (~(T1i2z4[9] & Hf5wx4));
assign Hf5wx4 = (~(Yz4wx4 & hwdata_o[9]));
assign Nevvx4 = (V15wx4 | Of5wx4);
assign Of5wx4 = (!hwdata_o[9]);
assign hwdata_o[9] = (Yd5wx4 ? Vf5wx4 : Htyvx4);
assign Ldvvx4 = (Uevvx4 | Vbovx4);
assign B0ivx4 = (Tavvx4 & Cg5wx4);
assign Cg5wx4 = (~(Jg5wx4 & Qg5wx4));
assign Qg5wx4 = (~(irq_i[10] & Mavvx4));
assign Mavvx4 = (!D3i2z4[10]);
assign Jg5wx4 = (Vbvvx4 & Xg5wx4);
assign Xg5wx4 = (~(T1i2z4[10] & Eh5wx4));
assign Eh5wx4 = (~(Yz4wx4 & hwdata_o[10]));
assign Vbvvx4 = (V15wx4 | Lh5wx4);
assign Lh5wx4 = (!hwdata_o[10]);
assign hwdata_o[10] = (Yd5wx4 ? Zh5wx4 : Sh5wx4);
assign Tavvx4 = (Ccvvx4 | Vbovx4);
assign Uzhvx4 = (B8vvx4 & Gi5wx4);
assign Gi5wx4 = (~(Ni5wx4 & Ui5wx4));
assign Ui5wx4 = (~(irq_i[11] & U7vvx4));
assign U7vvx4 = (!D3i2z4[11]);
assign Ni5wx4 = (D9vvx4 & Bj5wx4);
assign Bj5wx4 = (~(T1i2z4[11] & Ij5wx4));
assign Ij5wx4 = (~(Yz4wx4 & hwdata_o[11]));
assign D9vvx4 = (V15wx4 | Pj5wx4);
assign Pj5wx4 = (!hwdata_o[11]);
assign hwdata_o[11] = (Yd5wx4 ? Dk5wx4 : Wj5wx4);
assign B8vvx4 = (K9vvx4 | Vbovx4);
assign Nzhvx4 = (Lkvvx4 & Kk5wx4);
assign Kk5wx4 = (~(Rk5wx4 & Yk5wx4));
assign Yk5wx4 = (~(irq_i[12] & Ekvvx4));
assign Ekvvx4 = (!D3i2z4[12]);
assign Rk5wx4 = (Nlvvx4 & Fl5wx4);
assign Fl5wx4 = (~(T1i2z4[12] & Ml5wx4));
assign Ml5wx4 = (~(Yz4wx4 & hwdata_o[12]));
assign Nlvvx4 = (V15wx4 | Tl5wx4);
assign Tl5wx4 = (!hwdata_o[12]);
assign hwdata_o[12] = (Yd5wx4 ? Hm5wx4 : Am5wx4);
assign Lkvvx4 = (Ulvvx4 | Vbovx4);
assign Gzhvx4 = (P9uvx4 & Om5wx4);
assign Om5wx4 = (~(Vm5wx4 & Cn5wx4));
assign Cn5wx4 = (~(irq_i[13] & I9uvx4));
assign I9uvx4 = (!D3i2z4[13]);
assign Vm5wx4 = (Rauvx4 & Jn5wx4);
assign Jn5wx4 = (~(T1i2z4[13] & Qn5wx4));
assign Qn5wx4 = (~(Yz4wx4 & hwdata_o[13]));
assign Rauvx4 = (V15wx4 | Xn5wx4);
assign Xn5wx4 = (!hwdata_o[13]);
assign hwdata_o[13] = (Yd5wx4 ? Lo5wx4 : Eo5wx4);
assign P9uvx4 = (Yauvx4 | Vbovx4);
assign Zyhvx4 = (Awvvx4 & So5wx4);
assign So5wx4 = (~(Zo5wx4 & Gp5wx4));
assign Gp5wx4 = (~(irq_i[14] & Tvvvx4));
assign Tvvvx4 = (!D3i2z4[14]);
assign Zo5wx4 = (Cxvvx4 & Np5wx4);
assign Np5wx4 = (~(T1i2z4[14] & Up5wx4));
assign Up5wx4 = (~(Yz4wx4 & hwdata_o[14]));
assign hwdata_o[14] = (!Bq5wx4);
assign Cxvvx4 = (V15wx4 | Bq5wx4);
assign Bq5wx4 = (Iq5wx4 & Pq5wx4);
assign Iq5wx4 = (Wq5wx4 | S71wx4);
assign Awvvx4 = (Jxvvx4 | Vbovx4);
assign Syhvx4 = (Q6uvx4 & Dr5wx4);
assign Dr5wx4 = (~(Kr5wx4 & Rr5wx4));
assign Rr5wx4 = (~(irq_i[15] & J6uvx4));
assign J6uvx4 = (!D3i2z4[15]);
assign Kr5wx4 = (Z7uvx4 & Yr5wx4);
assign Yr5wx4 = (~(T1i2z4[15] & Fs5wx4));
assign Fs5wx4 = (~(Yz4wx4 & hwdata_o[15]));
assign Yz4wx4 = (Ms5wx4 & Ts5wx4);
assign Ms5wx4 = (~(Rgovx4 | Ctsvx4));
assign Z7uvx4 = (V15wx4 | At5wx4);
assign At5wx4 = (!hwdata_o[15]);
assign hwdata_o[15] = (Yd5wx4 ? Ot5wx4 : Ht5wx4);
assign V15wx4 = (!D9ovx4);
assign D9ovx4 = (Vt5wx4 & Ts5wx4);
assign Vt5wx4 = (~(Ctsvx4 | Xahvx4));
assign Ctsvx4 = (!Mf8vx4);
assign Q6uvx4 = (G8uvx4 | Vbovx4);
assign Vbovx4 = (~(Hg4wx4 & O4ovx4));
assign Hg4wx4 = (Cu5wx4 & Ju5wx4);
assign Cu5wx4 = (~(Tv2wx4 | Us2wx4));
assign Lyhvx4 = (!Qu5wx4);
assign Qu5wx4 = (Ccovx4 ? Ev5wx4 : Xu5wx4);
assign Xu5wx4 = (Lv5wx4 & Sv5wx4);
assign Sv5wx4 = (Zv5wx4 & Gw5wx4);
assign Gw5wx4 = (Nw5wx4 & Uw5wx4);
assign Uw5wx4 = (~(Bx5wx4 & Ix5wx4));
assign Bx5wx4 = (Px5wx4 & Wx5wx4);
assign Wx5wx4 = (R89vx4 ^ Dy5wx4);
assign Nw5wx4 = (~(Ky5wx4 | Ry5wx4));
assign Ky5wx4 = (!Yy5wx4);
assign Zv5wx4 = (Fz5wx4 & Mz5wx4);
assign Mz5wx4 = (~(Tz5wx4 & Liqvx4));
assign Tz5wx4 = (~(T93wx4 | U9gvx4));
assign Fz5wx4 = (A06wx4 & H06wx4);
assign H06wx4 = (~(O06wx4 & V06wx4));
assign O06wx4 = (Cf9vx4 & C16wx4);
assign C16wx4 = (J16wx4 | Qfsvx4);
assign A06wx4 = (~(Q16wx4 & X16wx4));
assign Q16wx4 = (E26wx4 & Xmsvx4);
assign E26wx4 = (V1yvx4 | L5wvx4);
assign Lv5wx4 = (L26wx4 & S26wx4);
assign S26wx4 = (Z26wx4 & G36wx4);
assign G36wx4 = (~(Sy2wx4 & N36wx4));
assign N36wx4 = (~(U36wx4 & B46wx4));
assign B46wx4 = (~(Liqvx4 & I46wx4));
assign I46wx4 = (~(Ujxvx4 & P46wx4));
assign P46wx4 = (Rexvx4 | Mj8vx4);
assign Z26wx4 = (W46wx4 & D56wx4);
assign D56wx4 = (~(Wdqvx4 & K56wx4));
assign K56wx4 = (~(R56wx4 & Y56wx4));
assign Y56wx4 = (~(F66wx4 & M66wx4));
assign F66wx4 = (P03wx4 & Hgxvx4);
assign R56wx4 = (Jppvx4 | Z6gvx4);
assign W46wx4 = (~(O9qvx4 & T66wx4));
assign T66wx4 = (~(A76wx4 & H76wx4));
assign H76wx4 = (~(O76wx4 & Eiqvx4));
assign L26wx4 = (V76wx4 & C86wx4);
assign C86wx4 = (~(Ilpvx4 & Jp3wx4));
assign Eyhvx4 = (J86wx4 & Q86wx4);
assign Q86wx4 = (~(X86wx4 & E96wx4));
assign E96wx4 = (L96wx4 & S96wx4);
assign S96wx4 = (Z96wx4 & Ga6wx4);
assign Ga6wx4 = (Fzyvx4 & Og4wx4);
assign Z96wx4 = (Na6wx4 & Ua6wx4);
assign Ua6wx4 = (~(Bb6wx4 & Ib6wx4));
assign Ib6wx4 = (~(Us2wx4 | Rexvx4));
assign Bb6wx4 = (~(Pxyvx4 | U0ovx4));
assign Na6wx4 = (~(Pb6wx4 & Q5gvx4));
assign Pb6wx4 = (T1xvx4 & M3ovx4);
assign L96wx4 = (Wb6wx4 & Dc6wx4);
assign Dc6wx4 = (~(Kc6wx4 & R7qvx4));
assign Kc6wx4 = (~(Rc6wx4 & Yc6wx4));
assign Yc6wx4 = (Fd6wx4 & Md6wx4);
assign Md6wx4 = (~(Td6wx4 & Bzwvx4));
assign Td6wx4 = (~(Zjwvx4 | Ho8vx4));
assign Fd6wx4 = (Ae6wx4 & Ffxvx4);
assign Ffxvx4 = (~(He6wx4 & C9yvx4));
assign He6wx4 = (Oe6wx4 & Zrvvx4);
assign Rc6wx4 = (Ve6wx4 & Cf6wx4);
assign Cf6wx4 = (~(B1vvx4 & Qp3wx4));
assign Ve6wx4 = (Jf6wx4 | Gcqvx4);
assign Wb6wx4 = (Qf6wx4 & Xf6wx4);
assign Xf6wx4 = (~(Ncqvx4 & Eg6wx4));
assign Eg6wx4 = (~(Lg6wx4 & Sg6wx4));
assign Sg6wx4 = (Pxyvx4 | Zg6wx4);
assign Qf6wx4 = (~(Gh6wx4 & Nh6wx4));
assign Nh6wx4 = (~(Uh6wx4 & Bi6wx4));
assign Bi6wx4 = (~(Ii6wx4 & Pi6wx4));
assign Pi6wx4 = (Wi6wx4 & Dj6wx4);
assign Ii6wx4 = (Kj6wx4 & Rj6wx4);
assign Kj6wx4 = (~(Yj6wx4 | Fk6wx4));
assign Uh6wx4 = (~(Nkpvx4 | Mk6wx4));
assign X86wx4 = (Tk6wx4 & Al6wx4);
assign Al6wx4 = (Hl6wx4 & Ol6wx4);
assign Hl6wx4 = (Vl6wx4 & Cm6wx4);
assign Cm6wx4 = (~(Y13wx4 & Jm6wx4));
assign Jm6wx4 = (~(Qm6wx4 & Xm6wx4));
assign Xm6wx4 = (~(Sjwvx4 & En6wx4));
assign En6wx4 = (~(Ln6wx4 & Sn6wx4));
assign Sn6wx4 = (~(Zn6wx4 | Cf9vx4));
assign Ln6wx4 = (Go6wx4 & Ix5wx4);
assign Go6wx4 = (Y99vx4 ? J16wx4 : R89vx4);
assign Qm6wx4 = (No6wx4 & Uo6wx4);
assign Uo6wx4 = (~(Mgwvx4 & Bp6wx4));
assign Bp6wx4 = (~(Dfpvx4 & Ip6wx4));
assign Ip6wx4 = (Qfsvx4 | Bisvx4);
assign No6wx4 = (~(Aj9vx4 & Pp6wx4));
assign Pp6wx4 = (~(Wp6wx4 & Dq6wx4));
assign Dq6wx4 = (~(Kq6wx4 & Xmsvx4));
assign Kq6wx4 = (~(Rq6wx4 & Yq6wx4));
assign Yq6wx4 = (Qfsvx4 ? Mr6wx4 : Fr6wx4);
assign Mr6wx4 = (!Tr6wx4);
assign Fr6wx4 = (~(As6wx4 & Hs6wx4));
assign Hs6wx4 = (Os6wx4 & Mc9vx4);
assign As6wx4 = (~(Vs6wx4 | J8svx4));
assign Rq6wx4 = (Kg9vx4 & Ct6wx4);
assign Wp6wx4 = (~(Jt6wx4 & Qt6wx4));
assign Qt6wx4 = (~(Y99vx4 ^ Xt6wx4));
assign Jt6wx4 = (~(Blwvx4 | Kg9vx4));
assign Vl6wx4 = (A8yvx4 | K7xvx4);
assign Tk6wx4 = (~(Eu6wx4 | Lu6wx4));
assign Lu6wx4 = (Sh9vx4 ? Zu6wx4 : Su6wx4);
assign Zu6wx4 = (~(F1xvx4 | Epxvx4));
assign F1xvx4 = (~(Gv6wx4 & D83wx4));
assign Gv6wx4 = (Howvx4 & Nv6wx4);
assign Eu6wx4 = (~(Uv6wx4 & Bw6wx4));
assign J86wx4 = (O8gvx4 | hready_i);
assign Xxhvx4 = (!Iw6wx4);
assign Iw6wx4 = (Ccovx4 ? Izwvx4 : Pw6wx4);
assign Pw6wx4 = (Ww6wx4 & Dx6wx4);
assign Dx6wx4 = (Kx6wx4 & Rx6wx4);
assign Rx6wx4 = (Yx6wx4 & Fy6wx4);
assign Fy6wx4 = (My6wx4 & Ty6wx4);
assign Ty6wx4 = (~(Az6wx4 & Hz6wx4));
assign Hz6wx4 = (Oz6wx4 & Pswvx4);
assign Oz6wx4 = (~(Blwvx4 | Dmgvx4));
assign Az6wx4 = (Vz6wx4 & Ukpvx4);
assign Vz6wx4 = (Xt6wx4 ^ Y99vx4);
assign Xt6wx4 = (~(C07wx4 & J07wx4));
assign J07wx4 = (Q07wx4 ^ X07wx4);
assign X07wx4 = (E17wx4 & L17wx4);
assign L17wx4 = (~(Jwpvx4 | Ix5wx4));
assign Jwpvx4 = (~(Xwpvx4 | Zxpvx4));
assign Xwpvx4 = (!vis_apsr_o[0]);
assign E17wx4 = (S17wx4 & Z17wx4);
assign Z17wx4 = (Ud9vx4 | G27wx4);
assign S17wx4 = (N27wx4 | U27wx4);
assign U27wx4 = (Phh2z4 ? Dmh2z4[31] : Zwcvx4);
assign N27wx4 = (~(B37wx4 & Zxpvx4));
assign Zxpvx4 = (~(I37wx4 & P37wx4));
assign I37wx4 = (W37wx4 & D47wx4);
assign D47wx4 = (~(K47wx4 & R47wx4));
assign R47wx4 = (~(S4xvx4 | W5yvx4));
assign K47wx4 = (~(Y47wx4 | F57wx4));
assign W37wx4 = (~(M57wx4 & Ucqvx4));
assign M57wx4 = (~(T57wx4 | Izwvx4));
assign B37wx4 = (Zwcvx4 | Dmh2z4[31]);
assign Zwcvx4 = (A67wx4 & Donvx4);
assign Donvx4 = (~(H67wx4 & O67wx4));
assign O67wx4 = (V67wx4 & C77wx4);
assign C77wx4 = (J77wx4 & Q77wx4);
assign Q77wx4 = (~(Ffqvx4 & X77wx4));
assign J77wx4 = (J43wx4 | F3ovx4);
assign V67wx4 = (E87wx4 & L87wx4);
assign L87wx4 = (Wt2wx4 | Fjgvx4);
assign E87wx4 = (S87wx4 | Bl3wx4);
assign H67wx4 = (Z87wx4 & G97wx4);
assign G97wx4 = (S4xvx4 ? U97wx4 : N97wx4);
assign U97wx4 = (Ba7wx4 & Ia7wx4);
assign Ia7wx4 = (Us2wx4 | Fjgvx4);
assign Ba7wx4 = (~(Pa7wx4 | Dbgvx4));
assign N97wx4 = (~(D83wx4 & Pcyvx4));
assign Z87wx4 = (Wa7wx4 & O8gvx4);
assign Wa7wx4 = (Nggvx4 ? Db7wx4 : Sznvx4);
assign Q07wx4 = (~(Kb7wx4 & Rb7wx4));
assign Rb7wx4 = (Qb3wx4 ? Yb7wx4 : Gd3wx4);
assign Yb7wx4 = (!vis_apsr_o[3]);
assign Gd3wx4 = (Ev5wx4 ? Y5zvx4 : Fc7wx4);
assign Kb7wx4 = (Mc7wx4 & Tc7wx4);
assign Mc7wx4 = (Uasvx4 | Ud9vx4);
assign C07wx4 = (Ad7wx4 & Hd7wx4);
assign Hd7wx4 = (Od7wx4 | Vd7wx4);
assign Vd7wx4 = (Zqpvx4 ? Dtpvx4 : vis_apsr_o[1]);
assign Zqpvx4 = (~(Ce7wx4 & P37wx4));
assign P37wx4 = (Je7wx4 & Qe7wx4);
assign Qe7wx4 = (~(Cn8vx4 & Xe7wx4));
assign Xe7wx4 = (~(Ef7wx4 & Lf7wx4));
assign Ef7wx4 = (~(Sf7wx4 & Hw2wx4));
assign Sf7wx4 = (~(Vdgvx4 | Whgvx4));
assign Je7wx4 = (Zf7wx4 & Gg7wx4);
assign Ce7wx4 = (Ng7wx4 & Ug7wx4);
assign Ug7wx4 = (~(Cn8vx4 & Bh7wx4));
assign Bh7wx4 = (~(Ih7wx4 & Ph7wx4));
assign Ng7wx4 = (~(Vdgvx4 & Wh7wx4));
assign Wh7wx4 = (~(Di7wx4 & Ki7wx4));
assign Ki7wx4 = (~(Ri7wx4 & Wkxvx4));
assign Di7wx4 = (Yi7wx4 & B03wx4);
assign Yi7wx4 = (~(Xx2wx4 & Fj7wx4));
assign Fj7wx4 = (M3ovx4 | Sy2wx4);
assign Dtpvx4 = (Ev5wx4 ? Gy9vx4 : Mj7wx4);
assign Mj7wx4 = (~(Tj7wx4 & Ak7wx4));
assign Ak7wx4 = (~(Hk7wx4 & Ok7wx4));
assign Hk7wx4 = (~(Vk7wx4 | R2ovx4));
assign R2ovx4 = (!vis_apsr_o[1]);
assign Tj7wx4 = (~(Cl7wx4 & Jl7wx4));
assign Jl7wx4 = (~(Ql7wx4 & Xl7wx4));
assign Xl7wx4 = (~(Em7wx4 & Lm7wx4));
assign Em7wx4 = (Sm7wx4 & Zm7wx4);
assign Sm7wx4 = (~(Gn7wx4 & Nn7wx4));
assign Nn7wx4 = (Db7wx4 | Fc7wx4);
assign Fc7wx4 = (Un7wx4 & Bo7wx4);
assign Bo7wx4 = (Io7wx4 & Po7wx4);
assign Po7wx4 = (~(Wo7wx4 & Dp7wx4));
assign Wo7wx4 = (~(Kp7wx4 & Rp7wx4));
assign Rp7wx4 = (~(Yp7wx4 & Fq7wx4));
assign Kp7wx4 = (~(Mq7wx4 & Tq7wx4));
assign Io7wx4 = (~(Ar7wx4 & Hr7wx4));
assign Un7wx4 = (Or7wx4 & Vr7wx4);
assign Vr7wx4 = (Cs7wx4 | Js7wx4);
assign Or7wx4 = (Qs7wx4 | Xs7wx4);
assign Gn7wx4 = (Et7wx4 | Mcgvx4);
assign Ql7wx4 = (Lt7wx4 | St7wx4);
assign St7wx4 = (Lm7wx4 & Zm7wx4);
assign Lm7wx4 = (~(Zt7wx4 & Gu7wx4));
assign Zt7wx4 = (!Vk7wx4);
assign Lt7wx4 = (F3ovx4 ? Et7wx4 : Nu7wx4);
assign Et7wx4 = (Uu7wx4 & Bv7wx4);
assign Bv7wx4 = (Iv7wx4 & Pv7wx4);
assign Pv7wx4 = (~(Wv7wx4 & Dw7wx4));
assign Wv7wx4 = (Yw7wx4 ? Rw7wx4 : Kw7wx4);
assign Iv7wx4 = (~(Fx7wx4 & Tq7wx4));
assign Uu7wx4 = (Mx7wx4 & Tx7wx4);
assign Tx7wx4 = (~(Ay7wx4 & Hy7wx4));
assign Mx7wx4 = (~(Oy7wx4 & Vy7wx4));
assign Oy7wx4 = (Fq7wx4 & Cz7wx4);
assign Nu7wx4 = (Jz7wx4 & Qz7wx4);
assign Qz7wx4 = (Xz7wx4 & E08wx4);
assign E08wx4 = (~(L08wx4 & Vy7wx4));
assign L08wx4 = (S08wx4 & Cz7wx4);
assign Xz7wx4 = (~(Ay7wx4 & Z08wx4));
assign Jz7wx4 = (G18wx4 & N18wx4);
assign N18wx4 = (~(Fx7wx4 & U18wx4));
assign G18wx4 = (~(Dw7wx4 & B28wx4));
assign Cl7wx4 = (Zm7wx4 | Vk7wx4);
assign Od7wx4 = (~(I28wx4 & Fdsvx4));
assign I28wx4 = (~(Fb9vx4 ^ Qfsvx4));
assign Ad7wx4 = (~(P28wx4 & W28wx4));
assign W28wx4 = (~(D38wx4 & Tc7wx4));
assign D38wx4 = (Qfsvx4 | Fb9vx4);
assign P28wx4 = (Hh3wx4 ^ K38wx4);
assign K38wx4 = (Qb3wx4 ? vis_apsr_o[2] : Ibzvx4);
assign Qb3wx4 = (R38wx4 & Op2wx4);
assign Op2wx4 = (~(Y38wx4 & Wkxvx4));
assign R38wx4 = (~(Cn8vx4 & F48wx4));
assign F48wx4 = (~(M48wx4 & T48wx4));
assign T48wx4 = (A58wx4 & H58wx4);
assign H58wx4 = (O58wx4 & B03wx4);
assign B03wx4 = (~(Z6gvx4 & U0ovx4));
assign A58wx4 = (V58wx4 & Lf7wx4);
assign Lf7wx4 = (~(C68wx4 & Z6gvx4));
assign C68wx4 = (J68wx4 & Q68wx4);
assign J68wx4 = (M93wx4 | S4xvx4);
assign V58wx4 = (Q68wx4 | S4xvx4);
assign M48wx4 = (X68wx4 & Ih7wx4);
assign Ih7wx4 = (E78wx4 | Whgvx4);
assign X68wx4 = (L78wx4 & S78wx4);
assign S78wx4 = (~(Xx2wx4 & W5yvx4));
assign L78wx4 = (~(Ucqvx4 & Hw2wx4));
assign Ibzvx4 = (!Z78wx4);
assign Z78wx4 = (Ev5wx4 ? N88wx4 : G88wx4);
assign N88wx4 = (~(U88wx4 & B98wx4));
assign B98wx4 = (I98wx4 & P98wx4);
assign P98wx4 = (W98wx4 & Da8wx4);
assign Da8wx4 = (Ka8wx4 & Ra8wx4);
assign Ra8wx4 = (~(Ya1wx4 | Xk1wx4));
assign Xk1wx4 = (Ya8wx4 & Axnvx4);
assign Axnvx4 = (!Qk1wx4);
assign Ya8wx4 = (I5bvx4 ? Mb8wx4 : Fb8wx4);
assign Ya1wx4 = (Tb8wx4 & Mwnvx4);
assign Tb8wx4 = (E8bvx4 ? Mb8wx4 : Fb8wx4);
assign Ka8wx4 = (Cs0wx4 & G11wx4);
assign G11wx4 = (~(Ac8wx4 & Rvnvx4));
assign Ac8wx4 = (Lcbvx4 ? Mb8wx4 : Fb8wx4);
assign Cs0wx4 = (~(Hc8wx4 & Dvnvx4));
assign Hc8wx4 = (Hfbvx4 ? Mb8wx4 : Fb8wx4);
assign W98wx4 = (Oc8wx4 & Vc8wx4);
assign Vc8wx4 = (Z80wx4 & Ri0wx4);
assign Ri0wx4 = (~(Cd8wx4 & Iunvx4));
assign Cd8wx4 = (Dibvx4 ? Mb8wx4 : Fb8wx4);
assign Z80wx4 = (~(Jd8wx4 & Utnvx4));
assign Jd8wx4 = (Zkbvx4 ? Mb8wx4 : Fb8wx4);
assign Oc8wx4 = (Luzvx4 & Qd8wx4);
assign Qd8wx4 = (~(Xd8wx4 & Ee8wx4));
assign Ee8wx4 = (~(Le8wx4 & Se8wx4));
assign Se8wx4 = (Ze8wx4 & Gf8wx4);
assign Gf8wx4 = (Nf8wx4 & Uf8wx4);
assign Uf8wx4 = (Bg8wx4 & O7zvx4);
assign Bg8wx4 = (~(Ig8wx4 | Pg8wx4));
assign Nf8wx4 = (~(Dk5wx4 | Wj5wx4));
assign Ze8wx4 = (Wg8wx4 & Dh8wx4);
assign Dh8wx4 = (Kh8wx4 & Ze1wx4);
assign Kh8wx4 = (~(Rd5wx4 | Kd5wx4));
assign Wg8wx4 = (~(Ot5wx4 | Lo5wx4));
assign Le8wx4 = (Rh8wx4 & Yh8wx4);
assign Yh8wx4 = (Fi8wx4 & Mi8wx4);
assign Mi8wx4 = (Ti8wx4 & Hk0wx4);
assign Ti8wx4 = (~(Aj8wx4 | Hj8wx4));
assign Fi8wx4 = (~(Oj8wx4 | Vj8wx4));
assign Oj8wx4 = (!W21wx4);
assign Rh8wx4 = (Ck8wx4 & Jk8wx4);
assign Jk8wx4 = (~(Qk8wx4 | Xk8wx4));
assign Ck8wx4 = (~(El8wx4 | Ll8wx4));
assign Luzvx4 = (~(Sl8wx4 & Fpnvx4));
assign Sl8wx4 = (O2bvx4 ? Mb8wx4 : Fb8wx4);
assign I98wx4 = (Zl8wx4 & Gm8wx4);
assign Gm8wx4 = (Nm8wx4 & Um8wx4);
assign Um8wx4 = (~(Uozvx4 | J61wx4));
assign J61wx4 = (Bn8wx4 & Fwnvx4);
assign Bn8wx4 = (P9bvx4 ? Mb8wx4 : Fb8wx4);
assign Uozvx4 = (In8wx4 & Zsnvx4);
assign In8wx4 = (Kmbvx4 ? Mb8wx4 : Fb8wx4);
assign Nm8wx4 = (Pn8wx4 & Wn8wx4);
assign Wn8wx4 = (~(Lhyvx4 & Do8wx4));
assign Do8wx4 = (~(Ko8wx4 & Ro8wx4));
assign Ro8wx4 = (Yo8wx4 & Fp8wx4);
assign Fp8wx4 = (Mp8wx4 & Tp8wx4);
assign Tp8wx4 = (~(Aq8wx4 | Dmh2z4[3]));
assign Aq8wx4 = (Dmh2z4[6] | Dmh2z4[8]);
assign Mp8wx4 = (~(Dmh2z4[26] | Dmh2z4[30]));
assign Yo8wx4 = (Hq8wx4 & Oq8wx4);
assign Oq8wx4 = (~(Vq8wx4 | Dmh2z4[21]));
assign Vq8wx4 = (Dmh2z4[22] | Dmh2z4[25]);
assign Hq8wx4 = (~(Dmh2z4[19] | Dmh2z4[20]));
assign Ko8wx4 = (Cr8wx4 & Jr8wx4);
assign Jr8wx4 = (Qr8wx4 & Xr8wx4);
assign Xr8wx4 = (~(Es8wx4 | Dmh2z4[16]));
assign Es8wx4 = (Dmh2z4[17] | Dmh2z4[18]);
assign Qr8wx4 = (~(Dmh2z4[14] | Dmh2z4[15]));
assign Cr8wx4 = (Ls8wx4 & Ss8wx4);
assign Ss8wx4 = (~(Dmh2z4[12] | Dmh2z4[13]));
assign Ls8wx4 = (~(Dmh2z4[0] | Dmh2z4[11]));
assign Pn8wx4 = (~(Zs8wx4 & Fb8wx4));
assign Zs8wx4 = (~(Gt8wx4 & Nt8wx4));
assign Nt8wx4 = (Ut8wx4 & Bu8wx4);
assign Bu8wx4 = (Iu8wx4 & Pu8wx4);
assign Pu8wx4 = (Y3bvx4 | F32wx4);
assign Iu8wx4 = (Abbvx4 | P82wx4);
assign Ut8wx4 = (Wu8wx4 & Dv8wx4);
assign Dv8wx4 = (Hlzvx4 | Vnbvx4);
assign Wu8wx4 = (Ojbvx4 | Lf0wx4);
assign Gt8wx4 = (Kv8wx4 & Rv8wx4);
assign Rv8wx4 = (T6bvx4 | Pg1wx4);
assign Kv8wx4 = (Yv8wx4 & Fw8wx4);
assign Fw8wx4 = (Sgbvx4 | Wo0wx4);
assign Yv8wx4 = (Wdbvx4 | Hy0wx4);
assign Zl8wx4 = (Mw8wx4 & Cgyvx4);
assign Cgyvx4 = (Tw8wx4 & Ax8wx4);
assign Ax8wx4 = (Hx8wx4 & Ox8wx4);
assign Ox8wx4 = (~(Xd8wx4 & Htyvx4));
assign Hx8wx4 = (Vx8wx4 & Cy8wx4);
assign Cy8wx4 = (~(Jy8wx4 & Qy8wx4));
assign Qy8wx4 = (~(Yryvx4 | Xy8wx4));
assign Jy8wx4 = (vis_control_o & Ez8wx4);
assign Vx8wx4 = (~(Dmh2z4[1] & Lhyvx4));
assign Tw8wx4 = (Lz8wx4 & Sz8wx4);
assign Sz8wx4 = (~(Zz8wx4 & vis_ipsr_o[1]));
assign Lz8wx4 = (Punvx4 ? N09wx4 : G09wx4);
assign N09wx4 = (Ihh2z4 ? Tkzvx4 : Olzvx4);
assign G09wx4 = (~(X8zvx4 & Ihh2z4));
assign Ihh2z4 = (~(U09wx4 ^ B19wx4));
assign U09wx4 = (~(I19wx4 & P19wx4));
assign P19wx4 = (~(W19wx4 & Htyvx4));
assign I19wx4 = (D29wx4 & K29wx4);
assign K29wx4 = (~(Ml9vx4 & R29wx4));
assign D29wx4 = (~(Uz8vx4 & Y29wx4));
assign Mw8wx4 = (F39wx4 & M39wx4);
assign M39wx4 = (~(T39wx4 & Mb8wx4));
assign T39wx4 = (~(A49wx4 & H49wx4));
assign H49wx4 = (O49wx4 & V49wx4);
assign V49wx4 = (C59wx4 & J59wx4);
assign J59wx4 = (~(Y3bvx4 & Ronvx4));
assign Ronvx4 = (!F32wx4);
assign C59wx4 = (~(Abbvx4 & Yvnvx4));
assign Yvnvx4 = (!P82wx4);
assign O49wx4 = (Q59wx4 & X59wx4);
assign X59wx4 = (~(Vnbvx4 & Ssnvx4));
assign Q59wx4 = (~(Ojbvx4 & Bunvx4));
assign A49wx4 = (E69wx4 & L69wx4);
assign L69wx4 = (~(T6bvx4 & Twnvx4));
assign E69wx4 = (S69wx4 & Z69wx4);
assign Z69wx4 = (~(Sgbvx4 & Wunvx4));
assign S69wx4 = (~(Wdbvx4 & Kvnvx4));
assign F39wx4 = (~(X8zvx4 & G79wx4));
assign G79wx4 = (~(N79wx4 & U79wx4));
assign U79wx4 = (B89wx4 & I89wx4);
assign I89wx4 = (P89wx4 & W89wx4);
assign W89wx4 = (D99wx4 & K99wx4);
assign K99wx4 = (~(Qk1wx4 & I5bvx4));
assign I5bvx4 = (~(R99wx4 ^ B19wx4));
assign R99wx4 = (~(Y99wx4 & Fa9wx4));
assign Fa9wx4 = (Ma9wx4 | Gm1wx4);
assign Y99wx4 = (Ta9wx4 & Ab9wx4);
assign Ta9wx4 = (~(Mc9vx4 & Y29wx4));
assign Qk1wx4 = (Hb9wx4 & Ob9wx4);
assign Ob9wx4 = (~(Vb9wx4 & Cc9wx4));
assign Cc9wx4 = (~(Jc9wx4 & Qc9wx4));
assign Qc9wx4 = (Xc9wx4 & Ed9wx4);
assign Ed9wx4 = (Ld9wx4 & Sd9wx4);
assign Sd9wx4 = (~(Zd9wx4 & vis_r14_o[11]));
assign Ld9wx4 = (Ge9wx4 & Ne9wx4);
assign Ne9wx4 = (~(Ue9wx4 & vis_psp_o[9]));
assign Ge9wx4 = (~(Bf9wx4 & vis_msp_o[9]));
assign Xc9wx4 = (If9wx4 & Pf9wx4);
assign Pf9wx4 = (~(Wf9wx4 & vis_r12_o[11]));
assign If9wx4 = (~(Dg9wx4 & vis_r11_o[11]));
assign Jc9wx4 = (Kg9wx4 & Rg9wx4);
assign Rg9wx4 = (Yg9wx4 & Fh9wx4);
assign Fh9wx4 = (~(Mh9wx4 & vis_r10_o[11]));
assign Yg9wx4 = (~(Th9wx4 & vis_r9_o[11]));
assign Kg9wx4 = (Ai9wx4 & Hi9wx4);
assign Hi9wx4 = (~(Oi9wx4 & vis_r8_o[11]));
assign Hb9wx4 = (Vi9wx4 & Cj9wx4);
assign Cj9wx4 = (~(Gcdvx4 & Jj9wx4));
assign Vi9wx4 = (~(Qj9wx4 & Rddvx4));
assign D99wx4 = (Xj9wx4 & Ek9wx4);
assign Ek9wx4 = (~(F32wx4 & Y3bvx4));
assign Y3bvx4 = (~(Lk9wx4 ^ B19wx4));
assign Lk9wx4 = (~(Sk9wx4 & Zk9wx4));
assign Zk9wx4 = (Gl9wx4 & Nl9wx4);
assign Nl9wx4 = (~(Gr9vx4 & Ul9wx4));
assign Gl9wx4 = (~(R89vx4 & Y29wx4));
assign Sk9wx4 = (Bm9wx4 & Im9wx4);
assign Im9wx4 = (G6wvx4 | Pm9wx4);
assign Bm9wx4 = (Ma9wx4 | P12wx4);
assign F32wx4 = (Wm9wx4 & Dn9wx4);
assign Dn9wx4 = (~(Vb9wx4 & Kn9wx4));
assign Kn9wx4 = (~(Rn9wx4 & Yn9wx4));
assign Yn9wx4 = (Fo9wx4 & Mo9wx4);
assign Mo9wx4 = (To9wx4 & Ap9wx4);
assign Ap9wx4 = (~(Zd9wx4 & vis_r14_o[8]));
assign To9wx4 = (Hp9wx4 & Op9wx4);
assign Op9wx4 = (~(Ue9wx4 & vis_psp_o[6]));
assign Hp9wx4 = (~(Bf9wx4 & vis_msp_o[6]));
assign Fo9wx4 = (Vp9wx4 & Cq9wx4);
assign Cq9wx4 = (~(Wf9wx4 & vis_r12_o[8]));
assign Vp9wx4 = (~(Dg9wx4 & vis_r11_o[8]));
assign Rn9wx4 = (Jq9wx4 & Qq9wx4);
assign Qq9wx4 = (Xq9wx4 & Er9wx4);
assign Er9wx4 = (~(Mh9wx4 & vis_r10_o[8]));
assign Xq9wx4 = (~(Th9wx4 & vis_r9_o[8]));
assign Jq9wx4 = (Lr9wx4 & Sr9wx4);
assign Sr9wx4 = (~(Oi9wx4 & vis_r8_o[8]));
assign Wm9wx4 = (Zr9wx4 & Gs9wx4);
assign Gs9wx4 = (~(C8dvx4 & Jj9wx4));
assign Zr9wx4 = (~(Qj9wx4 & M9dvx4));
assign Xj9wx4 = (~(P82wx4 & Abbvx4));
assign Abbvx4 = (~(Ns9wx4 ^ B19wx4));
assign Ns9wx4 = (~(Us9wx4 & Bt9wx4));
assign Bt9wx4 = (Ma9wx4 | Z62wx4);
assign Us9wx4 = (It9wx4 & Ab9wx4);
assign It9wx4 = (~(Yo9vx4 & Y29wx4));
assign P82wx4 = (Pt9wx4 & Wt9wx4);
assign Wt9wx4 = (~(Vb9wx4 & Du9wx4));
assign Du9wx4 = (~(Ku9wx4 & Ru9wx4));
assign Ru9wx4 = (Yu9wx4 & Fv9wx4);
assign Fv9wx4 = (Mv9wx4 & Tv9wx4);
assign Tv9wx4 = (~(Zd9wx4 & vis_r14_o[15]));
assign Mv9wx4 = (Aw9wx4 & Hw9wx4);
assign Hw9wx4 = (~(Ue9wx4 & vis_psp_o[13]));
assign Aw9wx4 = (~(Bf9wx4 & vis_msp_o[13]));
assign Yu9wx4 = (Ow9wx4 & Vw9wx4);
assign Vw9wx4 = (~(Wf9wx4 & vis_r12_o[15]));
assign Ow9wx4 = (~(Dg9wx4 & vis_r11_o[15]));
assign Ku9wx4 = (Cx9wx4 & Jx9wx4);
assign Jx9wx4 = (Qx9wx4 & Xx9wx4);
assign Xx9wx4 = (~(Mh9wx4 & vis_r10_o[15]));
assign Qx9wx4 = (~(Th9wx4 & vis_r9_o[15]));
assign Cx9wx4 = (Ey9wx4 & Ly9wx4);
assign Ly9wx4 = (~(Oi9wx4 & vis_r8_o[15]));
assign Pt9wx4 = (Sy9wx4 & Zy9wx4);
assign Zy9wx4 = (~(Yhdvx4 & Jj9wx4));
assign Sy9wx4 = (~(Qj9wx4 & Jjdvx4));
assign P89wx4 = (Gz9wx4 & Nz9wx4);
assign Nz9wx4 = (~(Q8zvx4 & Dih2z4));
assign Gz9wx4 = (~(Euzvx4 & O2bvx4));
assign O2bvx4 = (~(Uz9wx4 ^ B19wx4));
assign Uz9wx4 = (~(B0awx4 & I0awx4));
assign I0awx4 = (P0awx4 & W0awx4);
assign W0awx4 = (Xy8wx4 | D1awx4);
assign P0awx4 = (~(Y29wx4 & D69vx4));
assign B0awx4 = (K1awx4 & R1awx4);
assign R1awx4 = (~(Gr9vx4 & Y1awx4));
assign K1awx4 = (Ma9wx4 | Uvzvx4);
assign B89wx4 = (F2awx4 & M2awx4);
assign M2awx4 = (T2awx4 & A3awx4);
assign A3awx4 = (~(Hlzvx4 & Vnbvx4));
assign Vnbvx4 = (~(H3awx4 & O3awx4));
assign H3awx4 = (Djzvx4 ? C4awx4 : V3awx4);
assign T2awx4 = (~(Nozvx4 & Kmbvx4));
assign Kmbvx4 = (~(J4awx4 & O3awx4));
assign J4awx4 = (Kqzvx4 ? C4awx4 : V3awx4);
assign F2awx4 = (Q4awx4 & X4awx4);
assign X4awx4 = (~(N90wx4 & Zkbvx4));
assign Zkbvx4 = (~(E5awx4 ^ B19wx4));
assign E5awx4 = (~(L5awx4 & S5awx4));
assign S5awx4 = (Ud9vx4 ? G6awx4 : Z5awx4);
assign L5awx4 = (N6awx4 & Ab9wx4);
assign N6awx4 = (Ma9wx4 | Wa0wx4);
assign Q4awx4 = (~(Lf0wx4 & Ojbvx4));
assign Ojbvx4 = (~(U6awx4 ^ B19wx4));
assign U6awx4 = (~(B7awx4 & I7awx4));
assign I7awx4 = (Ma9wx4 | Ce0wx4);
assign B7awx4 = (P7awx4 & Ab9wx4);
assign P7awx4 = (~(Wv9vx4 & Y29wx4));
assign N79wx4 = (W7awx4 & D8awx4);
assign D8awx4 = (K8awx4 & R8awx4);
assign R8awx4 = (Y8awx4 & F9awx4);
assign F9awx4 = (~(Fj0wx4 & Dibvx4));
assign Dibvx4 = (~(M9awx4 ^ B19wx4));
assign M9awx4 = (~(T9awx4 & Aaawx4));
assign Aaawx4 = (Ma9wx4 | Hk0wx4);
assign T9awx4 = (Haawx4 & Ab9wx4);
assign Haawx4 = (~(Su9vx4 & Y29wx4));
assign Y8awx4 = (~(Wo0wx4 & Sgbvx4));
assign Sgbvx4 = (~(Oaawx4 ^ B19wx4));
assign Oaawx4 = (~(Vaawx4 & Cbawx4));
assign Cbawx4 = (Ma9wx4 | Nn0wx4);
assign Vaawx4 = (Jbawx4 & Ab9wx4);
assign Jbawx4 = (~(Ot9vx4 & Y29wx4));
assign K8awx4 = (Qbawx4 & Xbawx4);
assign Xbawx4 = (~(Qs0wx4 & Hfbvx4));
assign Hfbvx4 = (~(Ecawx4 ^ B19wx4));
assign Ecawx4 = (~(Lcawx4 & Scawx4));
assign Scawx4 = (Ma9wx4 | St0wx4);
assign Lcawx4 = (Zcawx4 & Ab9wx4);
assign Zcawx4 = (~(Ks9vx4 & Y29wx4));
assign Qbawx4 = (~(Hy0wx4 & Wdbvx4));
assign Wdbvx4 = (~(Gdawx4 ^ B19wx4));
assign Gdawx4 = (~(Ndawx4 & Udawx4));
assign Udawx4 = (Ma9wx4 | Yw0wx4);
assign Ndawx4 = (Beawx4 & Ab9wx4);
assign Beawx4 = (~(Y29wx4 & Gr9vx4));
assign W7awx4 = (Ieawx4 & Peawx4);
assign Peawx4 = (Weawx4 & Dfawx4);
assign Dfawx4 = (~(U11wx4 & Lcbvx4));
assign Lcbvx4 = (~(Kfawx4 ^ B19wx4));
assign Kfawx4 = (~(Rfawx4 & Yfawx4));
assign Yfawx4 = (Ma9wx4 | W21wx4);
assign Rfawx4 = (Fgawx4 & Ab9wx4);
assign Fgawx4 = (~(Cq9vx4 & Y29wx4));
assign Weawx4 = (~(C61wx4 & P9bvx4));
assign P9bvx4 = (~(Mgawx4 ^ B19wx4));
assign Mgawx4 = (~(Tgawx4 & Ahawx4));
assign Ahawx4 = (Ma9wx4 | S71wx4);
assign Tgawx4 = (Hhawx4 & Ab9wx4);
assign Hhawx4 = (~(Un9vx4 & Y29wx4));
assign Ieawx4 = (Ohawx4 & Vhawx4);
assign Vhawx4 = (~(Ra1wx4 & E8bvx4));
assign E8bvx4 = (~(Ciawx4 ^ B19wx4));
assign Ciawx4 = (~(Jiawx4 & Qiawx4));
assign Qiawx4 = (Ma9wx4 | Hc1wx4);
assign Jiawx4 = (Xiawx4 & Ab9wx4);
assign Xiawx4 = (~(Qm9vx4 & Y29wx4));
assign Ohawx4 = (~(Pg1wx4 & T6bvx4));
assign T6bvx4 = (~(Ejawx4 ^ B19wx4));
assign Ejawx4 = (~(Ljawx4 & Sjawx4));
assign Sjawx4 = (Ma9wx4 | Ze1wx4);
assign Ljawx4 = (Zjawx4 & Ab9wx4);
assign Zjawx4 = (~(Ml9vx4 & Y29wx4));
assign U88wx4 = (Gkawx4 & Nkawx4);
assign Nkawx4 = (Ukawx4 & Blawx4);
assign Blawx4 = (Ilawx4 & Plawx4);
assign Plawx4 = (Y5zvx4 & K5zvx4);
assign K5zvx4 = (Wlawx4 & Dmawx4);
assign Dmawx4 = (Kmawx4 & Rmawx4);
assign Rmawx4 = (~(Ymawx4 & vis_apsr_o[0]));
assign Kmawx4 = (Fnawx4 & Egzvx4);
assign Fnawx4 = (~(Dmh2z4[28] & Lhyvx4));
assign Wlawx4 = (Mnawx4 & Tnawx4);
assign Tnawx4 = (~(Xd8wx4 & Aoawx4));
assign Mnawx4 = (Esnvx4 ? Ooawx4 : Hoawx4);
assign Ooawx4 = (Whh2z4 ? Tkzvx4 : Olzvx4);
assign Hoawx4 = (~(X8zvx4 & Whh2z4));
assign Whh2z4 = (Aoawx4 ? Cpawx4 : Voawx4);
assign Y5zvx4 = (Jpawx4 & Qpawx4);
assign Qpawx4 = (Xpawx4 & Eqawx4);
assign Eqawx4 = (~(vis_apsr_o[3] & Ymawx4));
assign Xpawx4 = (Lqawx4 & Egzvx4);
assign Lqawx4 = (~(Dmh2z4[31] & Lhyvx4));
assign Jpawx4 = (Sqawx4 & Zqawx4);
assign Zqawx4 = (~(Xd8wx4 & Grawx4));
assign Sqawx4 = (A67wx4 ? Urawx4 : Nrawx4);
assign Urawx4 = (Phh2z4 ? Tkzvx4 : Olzvx4);
assign Nrawx4 = (~(X8zvx4 & Phh2z4));
assign Phh2z4 = (Grawx4 ? Cpawx4 : Voawx4);
assign Ilawx4 = (~(Giyvx4 | D5zvx4));
assign D5zvx4 = (~(Bsawx4 & Isawx4));
assign Isawx4 = (Psawx4 & Egzvx4);
assign Psawx4 = (~(Dmh2z4[7] & Lhyvx4));
assign Bsawx4 = (Wsawx4 & Dtawx4);
assign Dtawx4 = (~(Xd8wx4 & Ht5wx4));
assign Wsawx4 = (Yonvx4 ? Rtawx4 : Ktawx4);
assign Rtawx4 = (Ytawx4 & Fuawx4);
assign Ytawx4 = (Ugh2z4 ? Muawx4 : Alzvx4);
assign Ktawx4 = (~(X8zvx4 & Ugh2z4));
assign Ugh2z4 = (~(Tuawx4 ^ B19wx4));
assign Tuawx4 = (~(Avawx4 & Hvawx4));
assign Hvawx4 = (Ovawx4 & Vvawx4);
assign Vvawx4 = (Cwawx4 | D1awx4);
assign Ovawx4 = (~(Y29wx4 & K79vx4));
assign Avawx4 = (Jwawx4 & Qwawx4);
assign Qwawx4 = (~(Ks9vx4 & Y1awx4));
assign Y1awx4 = (!Xwawx4);
assign Jwawx4 = (~(W19wx4 & Ht5wx4));
assign Giyvx4 = (~(Exawx4 & Lxawx4));
assign Lxawx4 = (Sxawx4 & Egzvx4);
assign Sxawx4 = (~(Zxawx4 & Gyawx4));
assign Gyawx4 = (~(Xy8wx4 | Qm9vx4));
assign Zxawx4 = (Ez8wx4 & vis_primask_o);
assign Exawx4 = (Nyawx4 & Uyawx4);
assign Uyawx4 = (~(Zz8wx4 & vis_ipsr_o[0]));
assign Nyawx4 = (E1bvx4 ? Izawx4 : Bzawx4);
assign E1bvx4 = (Pzawx4 ^ Wzawx4);
assign Pzawx4 = (~(D0bwx4 & K0bwx4));
assign K0bwx4 = (~(Ik9vx4 & R29wx4));
assign D0bwx4 = (Ma9wx4 | Zhyvx4);
assign Izawx4 = (Oxnvx4 ? Tkzvx4 : Alzvx4);
assign Bzawx4 = (~(Fb8wx4 & Oxnvx4));
assign Ukawx4 = (R0bwx4 & Y0bwx4);
assign Y0bwx4 = (M50wx4 & L9zvx4);
assign L9zvx4 = (F1bwx4 & M1bwx4);
assign M1bwx4 = (~(vis_apsr_o[2] & Ymawx4));
assign F1bwx4 = (T1bwx4 & Egzvx4);
assign T1bwx4 = (~(A2bwx4 & Hqnvx4));
assign A2bwx4 = (Dih2z4 ? Mb8wx4 : Fb8wx4);
assign Dih2z4 = (H2bwx4 ? Cpawx4 : Voawx4);
assign M50wx4 = (O2bwx4 & V2bwx4);
assign V2bwx4 = (~(Zz8wx4 & vis_ipsr_o[3]));
assign O2bwx4 = (Sfh2z4 ? J3bwx4 : C3bwx4);
assign Sfh2z4 = (Q3bwx4 ^ Wzawx4);
assign Q3bwx4 = (~(X3bwx4 & E4bwx4));
assign E4bwx4 = (L4bwx4 & S4bwx4);
assign S4bwx4 = (~(Ml9vx4 & Z4bwx4));
assign L4bwx4 = (~(I29vx4 & Y29wx4));
assign X3bwx4 = (G5bwx4 & N5bwx4);
assign N5bwx4 = (U5bwx4 | Xwawx4);
assign G5bwx4 = (Ma9wx4 | R40wx4);
assign Ma9wx4 = (!W19wx4);
assign J3bwx4 = (Aqnvx4 ? Tkzvx4 : Alzvx4);
assign C3bwx4 = (~(Fb8wx4 & Aqnvx4));
assign Aqnvx4 = (~(B6bwx4 & I6bwx4));
assign I6bwx4 = (~(E1dvx4 & Jj9wx4));
assign B6bwx4 = (P6bwx4 & W6bwx4);
assign W6bwx4 = (~(Vb9wx4 & D7bwx4));
assign D7bwx4 = (~(K7bwx4 & R7bwx4));
assign R7bwx4 = (Y7bwx4 & F8bwx4);
assign F8bwx4 = (M8bwx4 & T8bwx4);
assign T8bwx4 = (~(vis_r14_o[3] & Zd9wx4));
assign M8bwx4 = (A9bwx4 & H9bwx4);
assign H9bwx4 = (~(vis_psp_o[1] & Ue9wx4));
assign A9bwx4 = (~(vis_msp_o[1] & Bf9wx4));
assign Y7bwx4 = (O9bwx4 & V9bwx4);
assign V9bwx4 = (~(vis_r12_o[3] & Wf9wx4));
assign O9bwx4 = (~(vis_r11_o[3] & Dg9wx4));
assign K7bwx4 = (Cabwx4 & Jabwx4);
assign Jabwx4 = (Qabwx4 & Xabwx4);
assign Xabwx4 = (~(vis_r10_o[3] & Mh9wx4));
assign Qabwx4 = (~(vis_r9_o[3] & Th9wx4));
assign Cabwx4 = (Ebbwx4 & Lbbwx4);
assign Lbbwx4 = (~(vis_r8_o[3] & Oi9wx4));
assign P6bwx4 = (~(O2dvx4 & Qj9wx4));
assign R0bwx4 = (Jr1wx4 & Xfzvx4);
assign Xfzvx4 = (Sbbwx4 & Zbbwx4);
assign Zbbwx4 = (Lsnvx4 ? Ncbwx4 : Gcbwx4);
assign Ncbwx4 = (Yih2z4 ? Tkzvx4 : Olzvx4);
assign Gcbwx4 = (~(X8zvx4 & Yih2z4));
assign Yih2z4 = (Ucbwx4 ? Cpawx4 : Voawx4);
assign Sbbwx4 = (Bdbwx4 & Idbwx4);
assign Idbwx4 = (~(Dmh2z4[27] & Lhyvx4));
assign Bdbwx4 = (Shyvx4 | Pdbwx4);
assign Jr1wx4 = (Wdbwx4 & Debwx4);
assign Debwx4 = (Kebwx4 & Rebwx4);
assign Rebwx4 = (~(Dmh2z4[2] & Lhyvx4));
assign Kebwx4 = (Yebwx4 & Ffbwx4);
assign Ffbwx4 = (~(Mfbwx4 & Tfbwx4));
assign Tfbwx4 = (O8gvx4 & Efgvx4);
assign Mfbwx4 = (Oy8vx4 & Agbwx4);
assign Yebwx4 = (~(Bpzvx4 & vis_control_o));
assign Wdbwx4 = (Hgbwx4 & Ogbwx4);
assign Ogbwx4 = (Qrnvx4 ? Chbwx4 : Vgbwx4);
assign Qrnvx4 = (~(Jhbwx4 & Qhbwx4));
assign Qhbwx4 = (~(Vb9wx4 & Xhbwx4));
assign Xhbwx4 = (~(Eibwx4 & Libwx4));
assign Libwx4 = (Sibwx4 & Zibwx4);
assign Zibwx4 = (Gjbwx4 & Njbwx4);
assign Njbwx4 = (~(vis_r14_o[2] & Zd9wx4));
assign Gjbwx4 = (Ujbwx4 & Bkbwx4);
assign Bkbwx4 = (~(vis_psp_o[0] & Ue9wx4));
assign Ujbwx4 = (~(vis_msp_o[0] & Bf9wx4));
assign Sibwx4 = (Ikbwx4 & Pkbwx4);
assign Pkbwx4 = (~(vis_r12_o[2] & Wf9wx4));
assign Ikbwx4 = (~(vis_r11_o[2] & Dg9wx4));
assign Eibwx4 = (Wkbwx4 & Dlbwx4);
assign Dlbwx4 = (Klbwx4 & Rlbwx4);
assign Rlbwx4 = (~(vis_r10_o[2] & Mh9wx4));
assign Klbwx4 = (~(vis_r9_o[2] & Th9wx4));
assign Wkbwx4 = (Ylbwx4 & Fmbwx4);
assign Fmbwx4 = (~(vis_r8_o[2] & Oi9wx4));
assign Jhbwx4 = (Mmbwx4 & Tmbwx4);
assign Tmbwx4 = (~(Uzcvx4 & Jj9wx4));
assign Mmbwx4 = (~(E1dvx4 & Qj9wx4));
assign Chbwx4 = (Anbwx4 & Fuawx4);
assign Anbwx4 = (Ngh2z4 ? Muawx4 : Alzvx4);
assign Vgbwx4 = (~(X8zvx4 & Ngh2z4));
assign Ngh2z4 = (~(Hnbwx4 ^ B19wx4));
assign Hnbwx4 = (~(Onbwx4 & Vnbwx4));
assign Vnbwx4 = (Cobwx4 & Jobwx4);
assign Jobwx4 = (~(Qm9vx4 & R29wx4));
assign R29wx4 = (~(Xwawx4 & Qobwx4));
assign Qobwx4 = (~(Xobwx4 & Epbwx4));
assign Epbwx4 = (Xx2wx4 & Dbgvx4);
assign Xobwx4 = (Ffqvx4 & O8gvx4);
assign Cobwx4 = (~(Ik9vx4 & Z4bwx4));
assign Onbwx4 = (Lpbwx4 & Spbwx4);
assign Spbwx4 = (~(B19vx4 & Y29wx4));
assign Lpbwx4 = (~(W19wx4 & Sh5wx4));
assign Hgbwx4 = (Zpbwx4 & Gqbwx4);
assign Gqbwx4 = (~(Xd8wx4 & Sh5wx4));
assign Zpbwx4 = (~(Zz8wx4 & vis_ipsr_o[2]));
assign Gkawx4 = (Nqbwx4 & Uqbwx4);
assign Uqbwx4 = (Brbwx4 & Irbwx4);
assign Irbwx4 = (Do1wx4 & Ox1wx4);
assign Ox1wx4 = (Prbwx4 & Wrbwx4);
assign Wrbwx4 = (Dsbwx4 & Egzvx4);
assign Dsbwx4 = (~(Dmh2z4[9] & Lhyvx4));
assign Prbwx4 = (Ksbwx4 & Rsbwx4);
assign Rsbwx4 = (~(Xd8wx4 & Vf5wx4));
assign Ksbwx4 = (Konvx4 ? Ftbwx4 : Ysbwx4);
assign Konvx4 = (~(Mtbwx4 & Ttbwx4));
assign Ttbwx4 = (~(M9dvx4 & Jj9wx4));
assign Mtbwx4 = (Aubwx4 & Hubwx4);
assign Hubwx4 = (~(Vb9wx4 & Oubwx4));
assign Oubwx4 = (~(Vubwx4 & Cvbwx4));
assign Cvbwx4 = (Jvbwx4 & Qvbwx4);
assign Qvbwx4 = (Xvbwx4 & Ewbwx4);
assign Ewbwx4 = (~(vis_r14_o[9] & Zd9wx4));
assign Xvbwx4 = (Lwbwx4 & Swbwx4);
assign Swbwx4 = (~(vis_psp_o[7] & Ue9wx4));
assign Lwbwx4 = (~(vis_msp_o[7] & Bf9wx4));
assign Jvbwx4 = (Zwbwx4 & Gxbwx4);
assign Gxbwx4 = (~(vis_r12_o[9] & Wf9wx4));
assign Zwbwx4 = (~(vis_r11_o[9] & Dg9wx4));
assign Vubwx4 = (Nxbwx4 & Uxbwx4);
assign Uxbwx4 = (Bybwx4 & Iybwx4);
assign Iybwx4 = (~(vis_r10_o[9] & Mh9wx4));
assign Bybwx4 = (~(vis_r9_o[9] & Th9wx4));
assign Nxbwx4 = (Pybwx4 & Wybwx4);
assign Wybwx4 = (~(vis_r8_o[9] & Oi9wx4));
assign Aubwx4 = (~(Wadvx4 & Qj9wx4));
assign Ftbwx4 = (Dzbwx4 & Fuawx4);
assign Dzbwx4 = (Bhh2z4 ? Muawx4 : Alzvx4);
assign Ysbwx4 = (~(X8zvx4 & Bhh2z4));
assign Bhh2z4 = (~(Kzbwx4 ^ B19wx4));
assign Kzbwx4 = (~(Rzbwx4 & Yzbwx4));
assign Yzbwx4 = (F0cwx4 & M0cwx4);
assign M0cwx4 = (~(Ks9vx4 & Ul9wx4));
assign Ul9wx4 = (!D1awx4);
assign F0cwx4 = (~(Y99vx4 & Y29wx4));
assign Rzbwx4 = (T0cwx4 & A1cwx4);
assign A1cwx4 = (~(Su9vx4 & H1cwx4));
assign T0cwx4 = (~(W19wx4 & Vf5wx4));
assign Do1wx4 = (O1cwx4 & V1cwx4);
assign V1cwx4 = (C2cwx4 & Egzvx4);
assign C2cwx4 = (~(Dmh2z4[10] & Lhyvx4));
assign O1cwx4 = (J2cwx4 & Q2cwx4);
assign Q2cwx4 = (~(Xd8wx4 & Zh5wx4));
assign J2cwx4 = (Hxnvx4 ? E3cwx4 : X2cwx4);
assign E3cwx4 = (L3cwx4 & Fuawx4);
assign L3cwx4 = (Mjh2z4 ? Muawx4 : Alzvx4);
assign X2cwx4 = (~(X8zvx4 & Mjh2z4));
assign Mjh2z4 = (~(S3cwx4 ^ B19wx4));
assign S3cwx4 = (~(Z3cwx4 & G4cwx4));
assign G4cwx4 = (~(W19wx4 & Zh5wx4));
assign Z3cwx4 = (N4cwx4 & U4cwx4);
assign U4cwx4 = (~(Fb9vx4 & Y29wx4));
assign N4cwx4 = (B5cwx4 | Pm9wx4);
assign Brbwx4 = (Yqzvx4 & Va3wx4);
assign Va3wx4 = (I5cwx4 & P5cwx4);
assign P5cwx4 = (W5cwx4 & Egzvx4);
assign W5cwx4 = (~(Dmh2z4[23] & Lhyvx4));
assign I5cwx4 = (D6cwx4 & K6cwx4);
assign K6cwx4 = (~(Xd8wx4 & R6cwx4));
assign D6cwx4 = (Ntnvx4 ? F7cwx4 : Y6cwx4);
assign F7cwx4 = (M7cwx4 & Fuawx4);
assign M7cwx4 = (Fjh2z4 ? Muawx4 : Alzvx4);
assign Y6cwx4 = (~(X8zvx4 & Fjh2z4));
assign Fjh2z4 = (~(T7cwx4 ^ B19wx4));
assign T7cwx4 = (~(A8cwx4 & H8cwx4));
assign H8cwx4 = (Dfpvx4 ? Z5awx4 : G6awx4);
assign Z5awx4 = (~(Y29wx4 & Dmwvx4));
assign A8cwx4 = (O8cwx4 & Ab9wx4);
assign O8cwx4 = (~(W19wx4 & R6cwx4));
assign Yqzvx4 = (V8cwx4 & C9cwx4);
assign C9cwx4 = (J9cwx4 & Egzvx4);
assign J9cwx4 = (~(Dmh2z4[24] & Lhyvx4));
assign V8cwx4 = (Q9cwx4 & X9cwx4);
assign X9cwx4 = (~(Xd8wx4 & Eacwx4));
assign Q9cwx4 = (Gtnvx4 ? Sacwx4 : Lacwx4);
assign Sacwx4 = (Zacwx4 & Fuawx4);
assign Zacwx4 = (Rih2z4 ? Muawx4 : Alzvx4);
assign Lacwx4 = (~(X8zvx4 & Rih2z4));
assign Rih2z4 = (Eacwx4 ? Cpawx4 : Voawx4);
assign Nqbwx4 = (Gbcwx4 & Fyzvx4);
assign Fyzvx4 = (Nbcwx4 & Ubcwx4);
assign Ubcwx4 = (Bccwx4 & Iccwx4);
assign Iccwx4 = (~(vis_ipsr_o[5] & Zz8wx4));
assign Bccwx4 = (Pccwx4 & Egzvx4);
assign Pccwx4 = (~(Dmh2z4[5] & Lhyvx4));
assign Nbcwx4 = (Wccwx4 & Ddcwx4);
assign Ddcwx4 = (~(Xd8wx4 & Eo5wx4));
assign Wccwx4 = (Mpnvx4 ? Rdcwx4 : Kdcwx4);
assign Rdcwx4 = (Zfh2z4 ? Tkzvx4 : Olzvx4);
assign Kdcwx4 = (~(X8zvx4 & Zfh2z4));
assign Zfh2z4 = (~(Ydcwx4 ^ B19wx4));
assign Ydcwx4 = (~(Fecwx4 & Mecwx4));
assign Mecwx4 = (Tecwx4 & Afcwx4);
assign Afcwx4 = (~(Un9vx4 & Z4bwx4));
assign Tecwx4 = (~(Y29wx4 & W49vx4));
assign Fecwx4 = (Hfcwx4 & Ofcwx4);
assign Ofcwx4 = (Cwawx4 | Xwawx4);
assign Hfcwx4 = (~(W19wx4 & Eo5wx4));
assign Gbcwx4 = (J00wx4 & Mdzvx4);
assign Mdzvx4 = (Vfcwx4 & Cgcwx4);
assign Cgcwx4 = (Jgcwx4 & Qgcwx4);
assign Qgcwx4 = (~(Ymawx4 & vis_apsr_o[1]));
assign Ymawx4 = (Ud3wx4 & Ez8wx4);
assign Ud3wx4 = (~(Qm9vx4 | Yo9vx4));
assign Jgcwx4 = (Xgcwx4 & Egzvx4);
assign Xgcwx4 = (~(Dmh2z4[29] & Lhyvx4));
assign Vfcwx4 = (Ehcwx4 & Lhcwx4);
assign Lhcwx4 = (~(Xd8wx4 & Shcwx4));
assign Ehcwx4 = (Xrnvx4 ? Gicwx4 : Zhcwx4);
assign Gicwx4 = (Nicwx4 & Fuawx4);
assign Nicwx4 = (Kih2z4 ? Muawx4 : Alzvx4);
assign Zhcwx4 = (~(X8zvx4 & Kih2z4));
assign Kih2z4 = (Shcwx4 ? Cpawx4 : Voawx4);
assign Cpawx4 = (~(O3awx4 & V3awx4));
assign V3awx4 = (~(W19wx4 & B19wx4));
assign Voawx4 = (~(O3awx4 & C4awx4));
assign O3awx4 = (Uicwx4 & Bjcwx4);
assign Bjcwx4 = (C4awx4 | W19wx4);
assign C4awx4 = (~(Ijcwx4 & Wzawx4));
assign Ijcwx4 = (G6awx4 & Ab9wx4);
assign Uicwx4 = (~(B19wx4 & Pjcwx4));
assign Pjcwx4 = (~(G6awx4 & Ab9wx4));
assign Ab9wx4 = (~(Bx9vx4 & H1cwx4));
assign H1cwx4 = (!Pm9wx4);
assign G6awx4 = (~(Bx9vx4 & Y29wx4));
assign J00wx4 = (Wjcwx4 & Dkcwx4);
assign Dkcwx4 = (Kkcwx4 & Rkcwx4);
assign Rkcwx4 = (~(Zz8wx4 & vis_ipsr_o[4]));
assign Zz8wx4 = (Ykcwx4 & Ez8wx4);
assign Ez8wx4 = (Flcwx4 & Mlcwx4);
assign Flcwx4 = (O8gvx4 & Tlcwx4);
assign Ykcwx4 = (~(Cppvx4 | Yo9vx4));
assign Kkcwx4 = (Amcwx4 & Egzvx4);
assign Egzvx4 = (!Bpzvx4);
assign Bpzvx4 = (Hmcwx4 & P03wx4);
assign Hmcwx4 = (O8gvx4 & Z6gvx4);
assign Amcwx4 = (~(Dmh2z4[4] & Lhyvx4));
assign Lhyvx4 = (~(Omcwx4 & Vmcwx4));
assign Vmcwx4 = (~(O8gvx4 & Cncwx4));
assign Cncwx4 = (Jncwx4 | Ps3wx4);
assign Jncwx4 = (S4xvx4 ? Qncwx4 : Auqvx4);
assign Qncwx4 = (~(Xncwx4 & Eocwx4));
assign Eocwx4 = (~(Locwx4 & F3ovx4));
assign Xncwx4 = (~(Socwx4 | Zocwx4));
assign Wjcwx4 = (Gpcwx4 & Npcwx4);
assign Npcwx4 = (~(Xd8wx4 & Am5wx4));
assign Xd8wx4 = (!Shyvx4);
assign Shyvx4 = (~(O8gvx4 & Upcwx4));
assign Upcwx4 = (~(Bqcwx4 & Iqcwx4));
assign Iqcwx4 = (~(Pcyvx4 & Nv6wx4));
assign Gpcwx4 = (Tpnvx4 ? Wqcwx4 : Pqcwx4);
assign Wqcwx4 = (Ggh2z4 ? Tkzvx4 : Olzvx4);
assign Tkzvx4 = (!Mb8wx4);
assign Mb8wx4 = (~(Fuawx4 & Muawx4));
assign Muawx4 = (Drcwx4 & Krcwx4);
assign Krcwx4 = (~(Rrcwx4 & Z6gvx4));
assign Rrcwx4 = (Yrcwx4 & B1ovx4);
assign Yrcwx4 = (U0ovx4 | Y38wx4);
assign Drcwx4 = (Fscwx4 | Lr2wx4);
assign Olzvx4 = (!Fb8wx4);
assign Fb8wx4 = (~(Fuawx4 & Alzvx4));
assign Alzvx4 = (!X8zvx4);
assign Fuawx4 = (Mscwx4 & Tscwx4);
assign Mscwx4 = (~(O8gvx4 & Atcwx4));
assign Atcwx4 = (~(Htcwx4 & Otcwx4));
assign Otcwx4 = (W5yvx4 ? Cucwx4 : Vtcwx4);
assign Cucwx4 = (~(Wkxvx4 & S4xvx4));
assign Vtcwx4 = (~(Pcyvx4 & Vdgvx4));
assign Htcwx4 = (Jucwx4 & Qucwx4);
assign Qucwx4 = (Jf6wx4 | O4ovx4);
assign Pqcwx4 = (~(X8zvx4 & Ggh2z4));
assign Ggh2z4 = (~(Xucwx4 ^ B19wx4));
assign B19wx4 = (!Wzawx4);
assign Wzawx4 = (O8gvx4 & Evcwx4);
assign Evcwx4 = (~(Lvcwx4 & Svcwx4));
assign Svcwx4 = (Zvcwx4 & Gwcwx4);
assign Gwcwx4 = (~(Nwcwx4 & Vdgvx4));
assign Nwcwx4 = (Uwcwx4 & U0ovx4);
assign Uwcwx4 = (~(Fscwx4 & Bxcwx4));
assign Bxcwx4 = (B1ovx4 | Nggvx4);
assign Zvcwx4 = (Ixcwx4 & H4ovx4);
assign H4ovx4 = (~(Pxcwx4 & Wxcwx4));
assign Ixcwx4 = (~(Dycwx4 & Zocwx4));
assign Dycwx4 = (Oe6wx4 & Cn8vx4);
assign Lvcwx4 = (T3ovx4 & Kycwx4);
assign Kycwx4 = (Jrnvx4 | Nggvx4);
assign T3ovx4 = (Rycwx4 & Yycwx4);
assign Yycwx4 = (~(X43wx4 & Kzxvx4));
assign Rycwx4 = (Fzcwx4 & Mzcwx4);
assign Mzcwx4 = (T57wx4 | Izwvx4);
assign Fzcwx4 = (~(Xx2wx4 & Hw2wx4));
assign Xucwx4 = (~(Tzcwx4 & A0dwx4));
assign A0dwx4 = (H0dwx4 & O0dwx4);
assign O0dwx4 = (~(Qm9vx4 & Z4bwx4));
assign Z4bwx4 = (~(D1awx4 & V0dwx4));
assign V0dwx4 = (~(O8gvx4 & C1dwx4));
assign C1dwx4 = (~(J1dwx4 & Q1dwx4));
assign Q1dwx4 = (X1dwx4 & E2dwx4);
assign E2dwx4 = (~(L2dwx4 & Whgvx4));
assign L2dwx4 = (S2dwx4 & Izwvx4);
assign S2dwx4 = (~(Z2dwx4 & G3dwx4));
assign G3dwx4 = (H33wx4 | W5yvx4);
assign X1dwx4 = (~(U9gvx4 & A2xvx4));
assign A2xvx4 = (B1vvx4 | Eiqvx4);
assign J1dwx4 = (N3dwx4 & U3dwx4);
assign U3dwx4 = (B4dwx4 | Wt2wx4);
assign N3dwx4 = (J43wx4 | Zrvvx4);
assign D1awx4 = (~(O8gvx4 & I4dwx4));
assign I4dwx4 = (~(P4dwx4 & W4dwx4));
assign W4dwx4 = (M3ovx4 ? K5dwx4 : D5dwx4);
assign K5dwx4 = (Lr2wx4 | Wt2wx4);
assign D5dwx4 = (~(R5dwx4 & D2ovx4));
assign P4dwx4 = (Y5dwx4 & F6dwx4);
assign F6dwx4 = (~(Bxyvx4 & Ucqvx4));
assign Bxyvx4 = (Mlcwx4 & Hw2wx4);
assign Mlcwx4 = (X77wx4 & Izwvx4);
assign Y5dwx4 = (~(Kzxvx4 & M6dwx4));
assign M6dwx4 = (T6dwx4 | R5dwx4);
assign T6dwx4 = (X43wx4 | Mcgvx4);
assign H0dwx4 = (~(P39vx4 & Y29wx4));
assign Y29wx4 = (A7dwx4 & H7dwx4);
assign H7dwx4 = (Hw2wx4 & F3ovx4);
assign A7dwx4 = (O8gvx4 & Vdgvx4);
assign Tzcwx4 = (O7dwx4 & V7dwx4);
assign V7dwx4 = (Xy8wx4 | Xwawx4);
assign Xwawx4 = (Pm9wx4 & C8dwx4);
assign C8dwx4 = (~(O8gvx4 & J8dwx4));
assign J8dwx4 = (~(Q8dwx4 & X8dwx4));
assign X8dwx4 = (~(E9dwx4 & Zrvvx4));
assign E9dwx4 = (~(L9dwx4 & S9dwx4));
assign S9dwx4 = (~(Z9dwx4 & W5yvx4));
assign Q8dwx4 = (Gadwx4 & Nadwx4);
assign Nadwx4 = (~(Hw2wx4 & Uadwx4));
assign Uadwx4 = (~(T57wx4 & Bbdwx4));
assign Bbdwx4 = (M3ovx4 | Nggvx4);
assign T57wx4 = (!Ibdwx4);
assign Gadwx4 = (~(Cn8vx4 & Pbdwx4));
assign Pbdwx4 = (~(Ph7wx4 & Wbdwx4));
assign Wbdwx4 = (B4dwx4 | Bl3wx4);
assign Pm9wx4 = (~(Dcdwx4 & O8gvx4));
assign Dcdwx4 = (~(N4yvx4 | Db7wx4));
assign O7dwx4 = (~(W19wx4 & Am5wx4));
assign W19wx4 = (O8gvx4 & Kcdwx4);
assign Kcdwx4 = (~(Rcdwx4 & Ycdwx4));
assign Ycdwx4 = (Fddwx4 & Mddwx4);
assign Mddwx4 = (~(Z6gvx4 & Tddwx4));
assign Tddwx4 = (~(Aedwx4 & Hedwx4));
assign Hedwx4 = (Fscwx4 | Oedwx4);
assign Aedwx4 = (Vedwx4 & Lr2wx4);
assign Lr2wx4 = (!Y38wx4);
assign Vedwx4 = (~(Mcgvx4 & Cfdwx4));
assign Cfdwx4 = (Us2wx4 | Vdgvx4);
assign Fddwx4 = (Jfdwx4 & Qfdwx4);
assign Qfdwx4 = (~(Xfdwx4 & Huqvx4));
assign Xfdwx4 = (~(Wt2wx4 | E78wx4));
assign Jfdwx4 = (~(Mcgvx4 & Egdwx4));
assign Egdwx4 = (~(F57wx4 & Lgdwx4));
assign Lgdwx4 = (~(D83wx4 & Q43wx4));
assign Rcdwx4 = (Sgdwx4 & Zgdwx4);
assign Zgdwx4 = (J43wx4 | Db7wx4);
assign Sgdwx4 = (S4xvx4 | Whgvx4);
assign X8zvx4 = (Ghdwx4 & Nhdwx4);
assign Nhdwx4 = (~(S4xvx4 | Whgvx4));
assign Ghdwx4 = (O8gvx4 & Qx2wx4);
assign G88wx4 = (~(Uhdwx4 & Bidwx4));
assign Bidwx4 = (Iidwx4 & Pidwx4);
assign Pidwx4 = (~(Widwx4 & Djdwx4));
assign Djdwx4 = (~(Kjdwx4 & Rjdwx4));
assign Rjdwx4 = (~(Yjdwx4 | Fkdwx4));
assign Yjdwx4 = (B28wx4 | Fq7wx4);
assign Kjdwx4 = (Mkdwx4 & Tkdwx4);
assign Mkdwx4 = (Oldwx4 ? Hldwx4 : Aldwx4);
assign Hldwx4 = (Vldwx4 & Cmdwx4);
assign Cmdwx4 = (~(Jmdwx4 | Rw7wx4));
assign Vldwx4 = (~(Qmdwx4 | Xmdwx4));
assign Aldwx4 = (Endwx4 & Lndwx4);
assign Lndwx4 = (~(Sndwx4 | Zndwx4));
assign Endwx4 = (~(Godwx4 | Nodwx4));
assign Widwx4 = (~(Uodwx4 & Bpdwx4));
assign Uodwx4 = (Ipdwx4 & Qs7wx4);
assign Iidwx4 = (Ppdwx4 & Wpdwx4);
assign Wpdwx4 = (~(Dqdwx4 & Kqdwx4));
assign Kqdwx4 = (~(Rqdwx4 & Yqdwx4));
assign Yqdwx4 = (~(Frdwx4 | Mrdwx4));
assign Frdwx4 = (U18wx4 | Hy7wx4);
assign Hy7wx4 = (!Xs7wx4);
assign Rqdwx4 = (Trdwx4 & Asdwx4);
assign Trdwx4 = (Oldwx4 ? Osdwx4 : Hsdwx4);
assign Osdwx4 = (Vsdwx4 & Ctdwx4);
assign Ctdwx4 = (~(Jtdwx4 | Qtdwx4));
assign Vsdwx4 = (~(Xtdwx4 | Eudwx4));
assign Hsdwx4 = (Ludwx4 & Sudwx4);
assign Sudwx4 = (~(Zudwx4 | Gvdwx4));
assign Ludwx4 = (~(Nvdwx4 | Uvdwx4));
assign Dqdwx4 = (~(Bwdwx4 & Iwdwx4));
assign Ppdwx4 = (~(Pwdwx4 & Wwdwx4));
assign Wwdwx4 = (~(Dxdwx4 & Kxdwx4));
assign Kxdwx4 = (~(Rxdwx4 | Yxdwx4));
assign Rxdwx4 = (S08wx4 | Tq7wx4);
assign Dxdwx4 = (Fydwx4 & Mydwx4);
assign Fydwx4 = (Oldwx4 ? Azdwx4 : Tydwx4);
assign Azdwx4 = (Hzdwx4 & Ozdwx4);
assign Ozdwx4 = (~(Vzdwx4 | Zndwx4));
assign Hzdwx4 = (~(C0ewx4 | Sndwx4));
assign Tydwx4 = (J0ewx4 & Q0ewx4);
assign Q0ewx4 = (~(Jtdwx4 | X0ewx4));
assign J0ewx4 = (~(E1ewx4 | Eudwx4));
assign Pwdwx4 = (~(Bwdwx4 & L1ewx4));
assign L1ewx4 = (S1ewx4 | Z1ewx4);
assign Uhdwx4 = (G2ewx4 & N2ewx4);
assign N2ewx4 = (~(U2ewx4 & B3ewx4));
assign B3ewx4 = (~(Cs7wx4 & I3ewx4));
assign G2ewx4 = (~(P3ewx4 & W3ewx4));
assign W3ewx4 = (~(D4ewx4 & K4ewx4));
assign K4ewx4 = (R4ewx4 & Y4ewx4);
assign Y4ewx4 = (~(F5ewx4 | M5ewx4));
assign R4ewx4 = (T5ewx4 & A6ewx4);
assign T5ewx4 = (~(H6ewx4 & O6ewx4));
assign O6ewx4 = (Kw7wx4 | Oldwx4);
assign D4ewx4 = (V6ewx4 & C7ewx4);
assign C7ewx4 = (~(J7ewx4 | Hr7wx4));
assign V6ewx4 = (Q7ewx4 & X7ewx4);
assign P3ewx4 = (~(E8ewx4 & L8ewx4));
assign L8ewx4 = (~(Ar7wx4 | Yp7wx4));
assign Ar7wx4 = (!S8ewx4);
assign E8ewx4 = (Z8ewx4 & S1ewx4);
assign My6wx4 = (~(G9ewx4 & N9ewx4));
assign G9ewx4 = (U9ewx4 & J8svx4);
assign U9ewx4 = (~(Baewx4 & Iaewx4));
assign Iaewx4 = (~(Paewx4 & Nywvx4));
assign Paewx4 = (~(Uasvx4 | Ud9vx4));
assign Baewx4 = (!Hh3wx4);
assign Yx6wx4 = (Waewx4 & Dbewx4);
assign Dbewx4 = (~(Kbewx4 & Ilpvx4));
assign Kbewx4 = (~(J43wx4 | B1ovx4));
assign Waewx4 = (~(Rbewx4 & Ih8vx4));
assign Rbewx4 = (~(Jppvx4 | Whgvx4));
assign Kx6wx4 = (Ybewx4 & Fcewx4);
assign Fcewx4 = (~(Mcewx4 & Tcewx4));
assign Tcewx4 = (~(Adewx4 & Hdewx4));
assign Hdewx4 = (Bl3wx4 ? Vdewx4 : Odewx4);
assign Vdewx4 = (Ceewx4 | Jeewx4);
assign Odewx4 = (~(Ucqvx4 & Efgvx4));
assign Adewx4 = (Qeewx4 & Xeewx4);
assign Xeewx4 = (Efewx4 | Nggvx4);
assign Qeewx4 = (F3ovx4 | Vdgvx4);
assign Ybewx4 = (Lfewx4 & Sfewx4);
assign Sfewx4 = (~(Px5wx4 & Zfewx4));
assign Zfewx4 = (~(Ggewx4 & Ngewx4));
assign Ngewx4 = (Zn6wx4 | Mc9vx4);
assign Ggewx4 = (Y99vx4 ? Fb9vx4 : Ugewx4);
assign Lfewx4 = (Bhewx4 | Ihewx4);
assign Ww6wx4 = (Phewx4 & Whewx4);
assign Whewx4 = (Diewx4 & Kiewx4);
assign Kiewx4 = (~(Soyvx4 & X16wx4));
assign Diewx4 = (Riewx4 & Yiewx4);
assign Yiewx4 = (~(Fjewx4 & Mjewx4));
assign Mjewx4 = (~(Tjewx4 & Akewx4));
assign Akewx4 = (F3ovx4 ? Okewx4 : Hkewx4);
assign Okewx4 = (~(Vkewx4 & R7qvx4));
assign Hkewx4 = (~(Clewx4 & Jlewx4));
assign Jlewx4 = (~(Efgvx4 & Qlewx4));
assign Qlewx4 = (~(Xlewx4 & Emewx4));
assign Tjewx4 = (Lmewx4 & Smewx4);
assign Smewx4 = (~(O76wx4 & B1vvx4));
assign Lmewx4 = (~(Zmewx4 & Bl3wx4));
assign Riewx4 = (~(Z9dwx4 & Gnewx4));
assign Phewx4 = (Nnewx4 & Unewx4);
assign Nnewx4 = (Boewx4 & Ioewx4);
assign Ioewx4 = (A76wx4 | Z6gvx4);
assign Boewx4 = (~(Huqvx4 & P6xvx4));
assign Qxhvx4 = (Poewx4 & Woewx4);
assign Woewx4 = (~(Dpewx4 & Kpewx4));
assign Kpewx4 = (Rpewx4 & Ypewx4);
assign Ypewx4 = (Fqewx4 & Mqewx4);
assign Mqewx4 = (Tqewx4 & Arewx4);
assign Tqewx4 = (~(Hrewx4 & A0zvx4));
assign Fqewx4 = (Orewx4 & Vrewx4);
assign Vrewx4 = (~(Csewx4 & Jsewx4));
assign Jsewx4 = (Aj9vx4 | Qsewx4);
assign Orewx4 = (~(Xsewx4 & Us2wx4));
assign Xsewx4 = (P6xvx4 | Liqvx4);
assign Rpewx4 = (Etewx4 & Ltewx4);
assign Ltewx4 = (Stewx4 & Ztewx4);
assign Ztewx4 = (~(Guewx4 & F3ovx4));
assign Guewx4 = (Howvx4 | Nuewx4);
assign Stewx4 = (~(Uuewx4 & Ud9vx4));
assign Etewx4 = (Bvewx4 & Ivewx4);
assign Ivewx4 = (Pvewx4 | Zg6wx4);
assign Bvewx4 = (~(Wvewx4 & Dwewx4));
assign Dwewx4 = (~(Kwewx4 & Rwewx4));
assign Rwewx4 = (Ywewx4 & Fxewx4);
assign Fxewx4 = (~(Sh9vx4 | R89vx4));
assign Ywewx4 = (~(Mxewx4 | Txewx4));
assign Mxewx4 = (Ud9vx4 & Vs6wx4);
assign Vs6wx4 = (~(Ayewx4 & Hyewx4));
assign Ayewx4 = (~(W49vx4 | K79vx4));
assign Kwewx4 = (Oyewx4 & G27wx4);
assign Oyewx4 = (~(Dfpvx4 | C1svx4));
assign Dpewx4 = (Vyewx4 & Czewx4);
assign Czewx4 = (Jzewx4 & Qzewx4);
assign Qzewx4 = (Xzewx4 & E0fwx4);
assign E0fwx4 = (~(Sh9vx4 & L0fwx4));
assign L0fwx4 = (~(S0fwx4 & Z0fwx4));
assign Z0fwx4 = (G1fwx4 & N1fwx4);
assign N1fwx4 = (~(U1fwx4 & Cn8vx4));
assign G1fwx4 = (~(Csewx4 & B2fwx4));
assign B2fwx4 = (~(I2fwx4 & P2fwx4));
assign P2fwx4 = (W2fwx4 & D3fwx4);
assign D3fwx4 = (~(K3fwx4 & Txewx4));
assign K3fwx4 = (~(Tc7wx4 | R89vx4));
assign W2fwx4 = (Ho3wx4 & Qfsvx4);
assign I2fwx4 = (R3fwx4 & Y3fwx4);
assign Y3fwx4 = (~(F4fwx4 & M4fwx4));
assign F4fwx4 = (~(J8svx4 | Fb9vx4));
assign S0fwx4 = (T4fwx4 & A5fwx4);
assign A5fwx4 = (Tc7wx4 | Icyvx4);
assign T4fwx4 = (~(G27wx4 & Xhxvx4));
assign Xzewx4 = (H5fwx4 | J8svx4);
assign Jzewx4 = (O5fwx4 & V5fwx4);
assign V5fwx4 = (~(T1xvx4 & Tlcwx4));
assign O5fwx4 = (Jf6wx4 | Msyvx4);
assign Vyewx4 = (C6fwx4 & J6fwx4);
assign J6fwx4 = (~(Q6fwx4 | X6fwx4));
assign X6fwx4 = (Ncqvx4 & Ju5wx4);
assign C6fwx4 = (~(E7fwx4 | L7fwx4));
assign L7fwx4 = (W5yvx4 ? Z7fwx4 : S7fwx4);
assign S7fwx4 = (Pcyvx4 & Socwx4);
assign E7fwx4 = (U0ovx4 ? Liqvx4 : G8fwx4);
assign G8fwx4 = (~(N8fwx4 & U8fwx4));
assign U8fwx4 = (B9fwx4 & I9fwx4);
assign I9fwx4 = (~(P9fwx4 & W9fwx4));
assign B9fwx4 = (Qhqvx4 | Hgxvx4);
assign N8fwx4 = (Dafwx4 & Kafwx4);
assign Kafwx4 = (~(Qp3wx4 & Sy2wx4));
assign Dafwx4 = (H33wx4 | Cn8vx4);
assign Poewx4 = (Whgvx4 | hready_i);
assign Jxhvx4 = (Yafwx4 ? Rafwx4 : Tjh2z4[3]);
assign Rafwx4 = (~(Fbfwx4 & Mbfwx4));
assign Mbfwx4 = (~(R89vx4 & Tbfwx4));
assign Tbfwx4 = (~(Acfwx4 & Hcfwx4));
assign Hcfwx4 = (Ocfwx4 | Fdsvx4);
assign Cxhvx4 = (~(Vcfwx4 & Cdfwx4));
assign Cdfwx4 = (Jdfwx4 & Qdfwx4);
assign Qdfwx4 = (~(Xdfwx4 & Dmh2z4[1]));
assign Jdfwx4 = (Eefwx4 & Lefwx4);
assign Eefwx4 = (Sefwx4 | C2rvx4);
assign C2rvx4 = (Zefwx4 & Gffwx4);
assign Gffwx4 = (Nffwx4 & Uffwx4);
assign Uffwx4 = (~(Bgfwx4 & Wjyvx4));
assign Nffwx4 = (Igfwx4 & Kkyvx4);
assign Igfwx4 = (~(Pgfwx4 & Ykyvx4));
assign Zefwx4 = (Wgfwx4 & Dhfwx4);
assign Dhfwx4 = (~(Khfwx4 & Omyvx4));
assign Wgfwx4 = (~(Rhfwx4 & Amyvx4));
assign Vcfwx4 = (Yhfwx4 & Fifwx4);
assign Fifwx4 = (~(Roh2z4[0] & Mifwx4));
assign Yhfwx4 = (Vlsvx4 | G6pvx4);
assign Vwhvx4 = (!Tifwx4);
assign Tifwx4 = (Ccovx4 ? W5yvx4 : Ajfwx4);
assign Ajfwx4 = (Hjfwx4 & Ojfwx4);
assign Ojfwx4 = (Vjfwx4 & Ckfwx4);
assign Ckfwx4 = (Jkfwx4 & Qkfwx4);
assign Qkfwx4 = (~(Vhpvx4 | Xkfwx4));
assign Jkfwx4 = (P7wvx4 & Elfwx4);
assign Vjfwx4 = (Llfwx4 & Slfwx4);
assign Slfwx4 = (~(Zlfwx4 & M1xvx4));
assign Zlfwx4 = (~(Gmfwx4 & Nmfwx4));
assign Nmfwx4 = (~(Umfwx4 & Ukpvx4));
assign Umfwx4 = (~(N4yvx4 | Mcgvx4));
assign Gmfwx4 = (~(Bnfwx4 & Nggvx4));
assign Llfwx4 = (Infwx4 & Pnfwx4);
assign Pnfwx4 = (~(Wnfwx4 & Clewx4));
assign Infwx4 = (~(B73wx4 & Dofwx4));
assign Dofwx4 = (~(Kofwx4 & Rofwx4));
assign Rofwx4 = (~(Yofwx4 & Qp3wx4));
assign Yofwx4 = (~(Fpfwx4 | Us2wx4));
assign Kofwx4 = (Jhxvx4 | J43wx4);
assign Hjfwx4 = (Mpfwx4 & Tpfwx4);
assign Tpfwx4 = (Aqfwx4 & Hqfwx4);
assign Hqfwx4 = (Oqfwx4 & Vqfwx4);
assign Vqfwx4 = (~(Whgvx4 & Crfwx4));
assign Crfwx4 = (~(Jrfwx4 & Qrfwx4));
assign Qrfwx4 = (~(Xrfwx4 & Ju5wx4));
assign Xrfwx4 = (~(Fjewx4 | U9gvx4));
assign Jrfwx4 = (Gjxvx4 | M3ovx4);
assign Oqfwx4 = (~(Bnfwx4 & Ucqvx4));
assign Aqfwx4 = (Esfwx4 & Lsfwx4);
assign Lsfwx4 = (~(C2yvx4 & Ssfwx4));
assign Ssfwx4 = (~(Zsfwx4 & Gtfwx4));
assign Gtfwx4 = (Ntfwx4 & Icyvx4);
assign Ntfwx4 = (~(Oowvx4 | Nkpvx4));
assign Zsfwx4 = (Utfwx4 & Bufwx4);
assign Bufwx4 = (Iufwx4 | Dfpvx4);
assign Utfwx4 = (Pufwx4 & Wufwx4);
assign Wufwx4 = (~(Dvfwx4 & Howvx4));
assign Dvfwx4 = (~(W5yvx4 | Aj9vx4));
assign Pufwx4 = (Kvfwx4 | Gwrvx4);
assign Esfwx4 = (~(Rvfwx4 & O4ovx4));
assign Rvfwx4 = (~(Yvfwx4 & Fwfwx4));
assign Fwfwx4 = (Mwfwx4 & Twfwx4);
assign Twfwx4 = (Axfwx4 & Hxfwx4);
assign Hxfwx4 = (~(Oxfwx4 & Rexvx4));
assign Oxfwx4 = (P9fwx4 & Ncqvx4);
assign Axfwx4 = (~(Cp3wx4 | Trsvx4));
assign Mwfwx4 = (Vxfwx4 & Cyfwx4);
assign Cyfwx4 = (~(Z7fwx4 & Jyfwx4));
assign Jyfwx4 = (~(Whgvx4 & Qyfwx4));
assign Qyfwx4 = (~(Ucqvx4 & Ujxvx4));
assign Vxfwx4 = (Xyfwx4 & Ezfwx4);
assign Ezfwx4 = (~(Lzfwx4 & U63wx4));
assign Lzfwx4 = (~(F3ovx4 | Cn8vx4));
assign Xyfwx4 = (~(Szfwx4 & Zzfwx4));
assign Szfwx4 = (~(Us2wx4 | Ki8vx4));
assign Yvfwx4 = (G0gwx4 & N0gwx4);
assign N0gwx4 = (U0gwx4 & B1gwx4);
assign B1gwx4 = (~(I1gwx4 & M1xvx4));
assign I1gwx4 = (~(P1gwx4 & W1gwx4));
assign W1gwx4 = (D2gwx4 & K2gwx4);
assign K2gwx4 = (~(Nkpvx4 & R2gwx4));
assign R2gwx4 = (~(Y2gwx4 & F3gwx4));
assign F3gwx4 = (M3gwx4 & T3gwx4);
assign T3gwx4 = (J8svx4 | Dj6wx4);
assign M3gwx4 = (~(A4gwx4 | H4gwx4));
assign Y2gwx4 = (O4gwx4 & V4gwx4);
assign V4gwx4 = (Y5svx4 | Fb9vx4);
assign O4gwx4 = (Mc9vx4 ? Ugewx4 : J16wx4);
assign D2gwx4 = (C5gwx4 & Avwvx4);
assign P1gwx4 = (J5gwx4 & Q5gwx4);
assign Q5gwx4 = (X5gwx4 | Ct6wx4);
assign J5gwx4 = (~(Hh3wx4 & Pyxvx4));
assign U0gwx4 = (E6gwx4 & L6gwx4);
assign L6gwx4 = (~(Pcyvx4 & S6gwx4));
assign S6gwx4 = (~(Ph7wx4 & Z6gwx4));
assign Z6gwx4 = (Oedwx4 | Sr2wx4);
assign E6gwx4 = (~(Howvx4 & G7gwx4));
assign G7gwx4 = (~(N7gwx4 & U7gwx4));
assign U7gwx4 = (B8gwx4 | Mcgvx4);
assign N7gwx4 = (I8gwx4 & Us2wx4);
assign I8gwx4 = (~(P8gwx4 & Rkgvx4));
assign P8gwx4 = (Vivvx4 & W5yvx4);
assign G0gwx4 = (W8gwx4 & D9gwx4);
assign D9gwx4 = (~(Wvewx4 & K9gwx4));
assign K9gwx4 = (~(R9gwx4 & Y9gwx4));
assign Y9gwx4 = (~(Cf9vx4 & Fagwx4));
assign Fagwx4 = (~(Magwx4 & Tagwx4));
assign Tagwx4 = (~(Abgwx4 ^ J8svx4));
assign Magwx4 = (Hbgwx4 & Obgwx4);
assign Obgwx4 = (Tc7wx4 | Qfsvx4);
assign Hbgwx4 = (J16wx4 | Mc9vx4);
assign R9gwx4 = (Vbgwx4 & Ccgwx4);
assign Ccgwx4 = (~(Jcgwx4 & Kg9vx4));
assign Jcgwx4 = (Y99vx4 & Qcgwx4);
assign Qcgwx4 = (~(Hyewx4 & Xcgwx4));
assign Xcgwx4 = (~(Edgwx4 & Ryrvx4));
assign Vbgwx4 = (~(Ldgwx4 & Qfsvx4));
assign Ldgwx4 = (~(Sdgwx4 & Fdsvx4));
assign Sdgwx4 = (~(Y5svx4 ^ Uasvx4));
assign W8gwx4 = (~(Pswvx4 & J8svx4));
assign Mpfwx4 = (Zdgwx4 & Nbyvx4);
assign Zdgwx4 = (Gegwx4 & Negwx4);
assign Negwx4 = (Z2zvx4 | Bswvx4);
assign Gegwx4 = (~(Wdqvx4 & Ju5wx4));
assign Owhvx4 = (!Uegwx4);
assign Uegwx4 = (Ccovx4 ? Us2wx4 : Bfgwx4);
assign Bfgwx4 = (Ifgwx4 & Pfgwx4);
assign Pfgwx4 = (Wfgwx4 & Dggwx4);
assign Dggwx4 = (Kggwx4 & Rggwx4);
assign Rggwx4 = (Yggwx4 & Fhgwx4);
assign Yggwx4 = (Vg4wx4 & Elfwx4);
assign Vg4wx4 = (~(M66wx4 & Wkxvx4));
assign Kggwx4 = (Mhgwx4 & Thgwx4);
assign Thgwx4 = (~(Aigwx4 & Higwx4));
assign Higwx4 = (~(Bdqvx4 | Ho8vx4));
assign Aigwx4 = (Oigwx4 & C2yvx4);
assign Mhgwx4 = (~(Vigwx4 & Cjgwx4));
assign Vigwx4 = (Jjgwx4 & Ukpvx4);
assign Wfgwx4 = (Qjgwx4 & Xjgwx4);
assign Xjgwx4 = (Ekgwx4 & Lkgwx4);
assign Lkgwx4 = (~(Skgwx4 & M66wx4));
assign Skgwx4 = (~(M3ovx4 | Nggvx4));
assign Ekgwx4 = (~(X16wx4 & Zkgwx4));
assign Zkgwx4 = (~(Avwvx4 & Glgwx4));
assign Glgwx4 = (~(Ud9vx4 & Nlgwx4));
assign Nlgwx4 = (~(Ulgwx4 & Bmgwx4));
assign Bmgwx4 = (~(Soyvx4 & Fb9vx4));
assign Avwvx4 = (~(Uuewx4 & Qfsvx4));
assign Qjgwx4 = (Imgwx4 & Pmgwx4);
assign Pmgwx4 = (~(Clewx4 & Wmgwx4));
assign Wmgwx4 = (Tlcwx4 | Dngwx4);
assign Dngwx4 = (Wdqvx4 & Kngwx4);
assign Imgwx4 = (~(Rngwx4 & Yngwx4));
assign Yngwx4 = (~(Fogwx4 & Mogwx4));
assign Mogwx4 = (~(Togwx4 & O4vvx4));
assign Togwx4 = (~(Apgwx4 & Hpgwx4));
assign Hpgwx4 = (Opgwx4 & Vpgwx4);
assign Opgwx4 = (~(Cqgwx4 & Howvx4));
assign Cqgwx4 = (Jqgwx4 & F3ovx4);
assign Jqgwx4 = (~(Qqgwx4 & Xqgwx4));
assign Xqgwx4 = (Xmsvx4 | Ho8vx4);
assign Apgwx4 = (Ergwx4 & Lrgwx4);
assign Lrgwx4 = (~(Q43wx4 & Dmgvx4));
assign Ergwx4 = (~(Pcyvx4 & W5yvx4));
assign Fogwx4 = (~(Srgwx4 & Gwrvx4));
assign Ifgwx4 = (Zrgwx4 & Gsgwx4);
assign Gsgwx4 = (Nsgwx4 & Usgwx4);
assign Usgwx4 = (Btgwx4 & Itgwx4);
assign Itgwx4 = (~(Ptgwx4 & Gnewx4));
assign Gnewx4 = (~(Jppvx4 & Wtgwx4));
assign Wtgwx4 = (~(Ilpvx4 & Z2zvx4));
assign Btgwx4 = (Dugwx4 & Kugwx4);
assign Kugwx4 = (~(O9qvx4 & Rugwx4));
assign Rugwx4 = (~(A76wx4 & Yugwx4));
assign Yugwx4 = (~(Fvgwx4 & C9yvx4));
assign Fvgwx4 = (~(Fscwx4 | Mvgwx4));
assign Dugwx4 = (Chxvx4 | Sznvx4);
assign Nsgwx4 = (Tvgwx4 & Awgwx4);
assign Awgwx4 = (~(Px5wx4 & Hwgwx4));
assign Hwgwx4 = (~(Owgwx4 & Vwgwx4));
assign Vwgwx4 = (~(Cxgwx4 & Ugewx4));
assign Cxgwx4 = (~(Ct6wx4 | Y99vx4));
assign Owgwx4 = (Jxgwx4 & Ho3wx4);
assign Ho3wx4 = (~(H4gwx4 & Fb9vx4));
assign Jxgwx4 = (!Qxgwx4);
assign Tvgwx4 = (~(Xxgwx4 & O4ovx4));
assign Xxgwx4 = (~(Eygwx4 & Lygwx4));
assign Lygwx4 = (Yyyvx4 & Sygwx4);
assign Eygwx4 = (Zygwx4 & Gzgwx4);
assign Gzgwx4 = (~(E44wx4 & A0zvx4));
assign Zygwx4 = (~(Nzgwx4 & Gh6wx4));
assign Zrgwx4 = (Uzgwx4 & B0hwx4);
assign B0hwx4 = (I0hwx4 & P0hwx4);
assign P0hwx4 = (~(Cf9vx4 & W0hwx4));
assign W0hwx4 = (~(D1hwx4 & K1hwx4));
assign K1hwx4 = (R1hwx4 & Y1hwx4);
assign Y1hwx4 = (~(F2hwx4 & M2hwx4));
assign M2hwx4 = (T2hwx4 & R7qvx4);
assign T2hwx4 = (~(A3hwx4 & H3hwx4));
assign H3hwx4 = (~(O3hwx4 & Fb9vx4));
assign A3hwx4 = (Ct6wx4 | J8svx4);
assign F2hwx4 = (Lxwvx4 & C2yvx4);
assign R1hwx4 = (~(V3hwx4 & Ihewx4));
assign Ihewx4 = (Edgwx4 & D69vx4);
assign Edgwx4 = (~(K79vx4 | R89vx4));
assign V3hwx4 = (~(Bhewx4 | Ryrvx4));
assign D1hwx4 = (C4hwx4 & J4hwx4);
assign J4hwx4 = (~(V06wx4 & Q4hwx4));
assign Q4hwx4 = (~(R89vx4 & X4hwx4));
assign X4hwx4 = (Qfsvx4 | N3svx4);
assign C4hwx4 = (~(X16wx4 & Ahwvx4));
assign I0hwx4 = (~(Pcyvx4 & E5hwx4));
assign E5hwx4 = (~(L5hwx4 & S5hwx4));
assign S5hwx4 = (Z5hwx4 & G6hwx4);
assign G6hwx4 = (~(R13wx4 & N6hwx4));
assign N6hwx4 = (Eznvx4 | U6hwx4);
assign Z5hwx4 = (B7hwx4 & I7hwx4);
assign I7hwx4 = (~(P7hwx4 & W7hwx4));
assign P7hwx4 = (D8hwx4 & K8hwx4);
assign B7hwx4 = (~(R8hwx4 & Sy2wx4));
assign R8hwx4 = (~(Bl3wx4 | Mj8vx4));
assign L5hwx4 = (Y8hwx4 & F9hwx4);
assign F9hwx4 = (~(Xhqvx4 & M9hwx4));
assign M9hwx4 = (~(Mv2wx4 & T9hwx4));
assign T9hwx4 = (~(Aahwx4 & W5yvx4));
assign Aahwx4 = (~(Vdgvx4 & Vivvx4));
assign Vivvx4 = (!C34wx4);
assign Y8hwx4 = (~(Hahwx4 & O4vvx4));
assign O4vvx4 = (!Rkgvx4);
assign Hahwx4 = (~(Oahwx4 & Vahwx4));
assign Vahwx4 = (~(Cbhwx4 & C2yvx4));
assign Cbhwx4 = (~(S4xvx4 | Z6gvx4));
assign Oahwx4 = (~(B73wx4 & O9qvx4));
assign Uzgwx4 = (~(Jbhwx4 | Qbhwx4));
assign Qbhwx4 = (~(S87wx4 | Pxyvx4));
assign Jbhwx4 = (U0ovx4 ? P5yvx4 : Xbhwx4);
assign Xbhwx4 = (~(Echwx4 & Lchwx4));
assign Lchwx4 = (~(Sy2wx4 & Kzxvx4));
assign Echwx4 = (Schwx4 & Zchwx4);
assign Zchwx4 = (Sznvx4 | B4dwx4);
assign Schwx4 = (~(Zmewx4 & Ujxvx4));
assign Hwhvx4 = (!Gdhwx4);
assign Gdhwx4 = (Ccovx4 ? M3ovx4 : Ndhwx4);
assign Ndhwx4 = (Udhwx4 & Behwx4);
assign Behwx4 = (Iehwx4 & Pehwx4);
assign Pehwx4 = (Wehwx4 & Dfhwx4);
assign Dfhwx4 = (~(Kfhwx4 & Rfhwx4));
assign Rfhwx4 = (Bnfwx4 | Yfhwx4);
assign Yfhwx4 = (Ilpvx4 & Us2wx4);
assign Kfhwx4 = (~(Dbgvx4 | Z6gvx4));
assign Wehwx4 = (~(Fghwx4 | B4zvx4));
assign B4zvx4 = (~(Pxyvx4 | M3ovx4));
assign Fghwx4 = (Mghwx4 & Emewx4);
assign Mghwx4 = (~(Zq3wx4 | S87wx4));
assign Iehwx4 = (Tghwx4 & Ahhwx4);
assign Ahhwx4 = (~(Hhhwx4 & Clewx4));
assign Hhhwx4 = (Xx2wx4 & Kngwx4);
assign Tghwx4 = (~(Ju5wx4 & Ohhwx4));
assign Ohhwx4 = (~(S4xvx4 & Vhhwx4));
assign Vhhwx4 = (Cihwx4 | Efgvx4);
assign Udhwx4 = (Jihwx4 & Qihwx4);
assign Qihwx4 = (Xihwx4 & Ejhwx4);
assign Ejhwx4 = (Vpgwx4 | U4yvx4);
assign Vpgwx4 = (~(Ljhwx4 & Dmgvx4));
assign Ljhwx4 = (~(U0ovx4 | Mcgvx4));
assign Xihwx4 = (Sjhwx4 & Zjhwx4);
assign Zjhwx4 = (~(Bnfwx4 & D2ovx4));
assign Bnfwx4 = (Pcyvx4 & Rngwx4);
assign Sjhwx4 = (~(Gkhwx4 & W5yvx4));
assign Gkhwx4 = (~(Nkhwx4 & Ukhwx4));
assign Ukhwx4 = (~(Blhwx4 & P6xvx4));
assign Blhwx4 = (~(Ilhwx4 | Efgvx4));
assign Nkhwx4 = (Plhwx4 & Agxvx4);
assign Plhwx4 = (~(Wlhwx4 & P9fwx4));
assign Jihwx4 = (Dmhwx4 & Kmhwx4);
assign Kmhwx4 = (Agxvx4 | Hgxvx4);
assign Agxvx4 = (~(Huqvx4 & Fjgvx4));
assign Dmhwx4 = (~(Rmhwx4 & O4ovx4));
assign Rmhwx4 = (~(Ymhwx4 & Fnhwx4));
assign Fnhwx4 = (Mnhwx4 & Tnhwx4);
assign Tnhwx4 = (Aohwx4 & Hohwx4);
assign Aohwx4 = (C5gwx4 & Oohwx4);
assign C5gwx4 = (~(Qoxvx4 & Lcpvx4));
assign Qoxvx4 = (~(Iufwx4 | Qfsvx4));
assign Mnhwx4 = (Vohwx4 & Cphwx4);
assign Cphwx4 = (~(Jphwx4 & Pcyvx4));
assign Jphwx4 = (U9gvx4 & Qphwx4);
assign Qphwx4 = (B1ovx4 | Tlcwx4);
assign Vohwx4 = (Xphwx4 & Eqhwx4);
assign Xphwx4 = (~(Lqhwx4 & Sqhwx4));
assign Sqhwx4 = (Qp3wx4 & O9qvx4);
assign Lqhwx4 = (~(Ujxvx4 | Fscwx4));
assign Ymhwx4 = (Zqhwx4 & Grhwx4);
assign Grhwx4 = (Nrhwx4 & Urhwx4);
assign Urhwx4 = (Jf6wx4 | Hq1wx4);
assign Nrhwx4 = (Bshwx4 & Ishwx4);
assign Ishwx4 = (~(Pshwx4 & Wshwx4));
assign Pshwx4 = (~(J8svx4 | Mc9vx4));
assign Bshwx4 = (Dthwx4 | Iufwx4);
assign Zqhwx4 = (~(Kthwx4 | Rthwx4));
assign Rthwx4 = (Qfsvx4 ? Pyxvx4 : Ythwx4);
assign Ythwx4 = (~(Tc7wx4 | Yj6wx4));
assign Kthwx4 = (~(Fuhwx4 & Muhwx4));
assign Muhwx4 = (~(A0zvx4 & Wdxvx4));
assign Fuhwx4 = (Izwvx4 ? Avhwx4 : Tuhwx4);
assign Avhwx4 = (Hvhwx4 & Ovhwx4);
assign Ovhwx4 = (~(Vvhwx4 & Fjewx4));
assign Vvhwx4 = (~(Oedwx4 | Fpfwx4));
assign Hvhwx4 = (~(U6hwx4 & Xx2wx4));
assign Tuhwx4 = (Cwhwx4 & Jwhwx4);
assign Jwhwx4 = (Qwhwx4 & Xwhwx4);
assign Xwhwx4 = (~(Ho8vx4 | Dmgvx4));
assign Qwhwx4 = (Exhwx4 & Lxhwx4);
assign Lxhwx4 = (~(Sxhwx4 & Fb9vx4));
assign Sxhwx4 = (Y5svx4 ? Gyhwx4 : Zxhwx4);
assign Gyhwx4 = (~(Bisvx4 | K79vx4));
assign Zxhwx4 = (~(Nyhwx4 & Uyhwx4));
assign Uyhwx4 = (B8gwx4 | N3svx4);
assign Nyhwx4 = (Dfpvx4 | Qfsvx4);
assign Exhwx4 = (~(Qsewx4 & Bzhwx4));
assign Bzhwx4 = (~(Izhwx4 & Rj6wx4));
assign Rj6wx4 = (~(C1svx4 ^ N3svx4));
assign Izhwx4 = (~(Fk6wx4 | Uasvx4));
assign Cwhwx4 = (Pzhwx4 & Wzhwx4);
assign Wzhwx4 = (Abgwx4 | Bisvx4);
assign Pzhwx4 = (D0iwx4 & K0iwx4);
assign K0iwx4 = (~(R0iwx4 & Lcpvx4));
assign R0iwx4 = (~(Y0iwx4 & F1iwx4));
assign F1iwx4 = (Kg9vx4 ? Bisvx4 : Lqwvx4);
assign Y0iwx4 = (M1iwx4 & T1iwx4);
assign T1iwx4 = (~(Oigwx4 & Fk6wx4));
assign M1iwx4 = (Ct6wx4 | Xmsvx4);
assign D0iwx4 = (~(Oigwx4 & Xmsvx4));
assign Awhvx4 = (Yafwx4 ? A2iwx4 : Tjh2z4[0]);
assign A2iwx4 = (~(H2iwx4 & O2iwx4));
assign O2iwx4 = (V2iwx4 & C3iwx4);
assign C3iwx4 = (J8svx4 | J3iwx4);
assign V2iwx4 = (~(Q3iwx4 & P39vx4));
assign H2iwx4 = (Fbfwx4 & X3iwx4);
assign X3iwx4 = (~(Uz8vx4 & E4iwx4));
assign Tvhvx4 = (~(L4iwx4 & S4iwx4));
assign S4iwx4 = (Z4iwx4 & G5iwx4);
assign G5iwx4 = (~(Xdfwx4 & Dmh2z4[30]));
assign Z4iwx4 = (N5iwx4 & Lefwx4);
assign N5iwx4 = (Sefwx4 | E9zvx4);
assign E9zvx4 = (U5iwx4 & B6iwx4);
assign B6iwx4 = (I6iwx4 & P6iwx4);
assign P6iwx4 = (~(W6iwx4 & D7iwx4));
assign I6iwx4 = (K7iwx4 & R7iwx4);
assign K7iwx4 = (~(Y7iwx4 & F8iwx4));
assign U5iwx4 = (M8iwx4 & T8iwx4);
assign T8iwx4 = (~(A9iwx4 & H9iwx4));
assign M8iwx4 = (~(O9iwx4 & V9iwx4));
assign L4iwx4 = (Caiwx4 & Jaiwx4);
assign Jaiwx4 = (~(Roh2z4[29] & Mifwx4));
assign Caiwx4 = (~(vis_pc_o[29] & Qaiwx4));
assign Mvhvx4 = (Xaiwx4 | Ebiwx4);
assign Ebiwx4 = (~(Lbiwx4 | Nggvx4));
assign Xaiwx4 = (Ccovx4 ? Dbgvx4 : Sbiwx4);
assign Sbiwx4 = (~(Zbiwx4 & Gciwx4));
assign Gciwx4 = (Nciwx4 & Uciwx4);
assign Uciwx4 = (Bdiwx4 & Idiwx4);
assign Idiwx4 = (~(Pdiwx4 & F3ovx4));
assign Pdiwx4 = (~(Elfwx4 & Wdiwx4));
assign Wdiwx4 = (~(Deiwx4 & Mcewx4));
assign Deiwx4 = (~(J43wx4 | Efgvx4));
assign Elfwx4 = (~(Howvx4 & B73wx4));
assign Bdiwx4 = (~(Keiwx4 & Cjgwx4));
assign Nciwx4 = (Reiwx4 & Yeiwx4);
assign Yeiwx4 = (~(Ffiwx4 & R7qvx4));
assign Ffiwx4 = (~(Mfiwx4 & Tfiwx4));
assign Tfiwx4 = (P7wvx4 | Qfsvx4);
assign Mfiwx4 = (Agiwx4 & Hgiwx4);
assign Hgiwx4 = (~(U1fwx4 & Ohwvx4));
assign Agiwx4 = (~(Vkewx4 & D2ovx4));
assign D2ovx4 = (O9qvx4 & Nggvx4);
assign Vkewx4 = (Ogiwx4 & Clewx4);
assign Ogiwx4 = (~(S87wx4 | Bl3wx4));
assign Reiwx4 = (~(Vgiwx4 & O4ovx4));
assign Vgiwx4 = (~(Chiwx4 & Jhiwx4));
assign Jhiwx4 = (Qhiwx4 & Yyyvx4);
assign Yyyvx4 = (Kvfwx4 | Nggvx4);
assign Qhiwx4 = (Hohwx4 & Xhiwx4);
assign Hohwx4 = (~(Eiiwx4 & Liiwx4));
assign Eiiwx4 = (~(Bqcwx4 | Msyvx4));
assign Chiwx4 = (Siiwx4 & Ziiwx4);
assign Ziiwx4 = (Kvfwx4 | Mv2wx4);
assign Siiwx4 = (Gjiwx4 & Mn3wx4);
assign Gjiwx4 = (~(A0zvx4 & Njiwx4));
assign Njiwx4 = (U63wx4 | Ujiwx4);
assign Zbiwx4 = (Bkiwx4 & Ikiwx4);
assign Ikiwx4 = (Pkiwx4 & Wkiwx4);
assign Wkiwx4 = (~(Qaqvx4 & Dliwx4));
assign Dliwx4 = (~(Kliwx4 & Rliwx4));
assign Rliwx4 = (Yliwx4 & Fmiwx4);
assign Fmiwx4 = (~(Ud9vx4 & Mmiwx4));
assign Mmiwx4 = (Tmiwx4 | Aniwx4);
assign Aniwx4 = (Fdsvx4 ? Wvewx4 : Hniwx4);
assign Hniwx4 = (~(B8gwx4 | Izwvx4));
assign Tmiwx4 = (~(Oniwx4 & Vniwx4));
assign Vniwx4 = (~(Coiwx4 & Q4wvx4));
assign Coiwx4 = (~(Ho8vx4 | Fb9vx4));
assign Oniwx4 = (Ulgwx4 | Dfpvx4);
assign Yliwx4 = (Joiwx4 & Qoiwx4);
assign Joiwx4 = (~(Xoiwx4 & Wvewx4));
assign Xoiwx4 = (~(Kg9vx4 | Y99vx4));
assign Kliwx4 = (~(Epiwx4 | Lpiwx4));
assign Lpiwx4 = (Xmsvx4 ? Oowvx4 : Spiwx4);
assign Spiwx4 = (Zpiwx4 & Csewx4);
assign Zpiwx4 = (Gqiwx4 & M1xvx4);
assign Gqiwx4 = (~(Nqiwx4 & Oigwx4));
assign Nqiwx4 = (Uqiwx4 & Briwx4);
assign Briwx4 = (~(Iriwx4 & Dj6wx4));
assign Iriwx4 = (~(Y5svx4 | Dy5wx4));
assign Dy5wx4 = (~(J8svx4 | K79vx4));
assign Uqiwx4 = (~(Y99vx4 & Priwx4));
assign Priwx4 = (~(Wriwx4 & Dsiwx4));
assign Dsiwx4 = (~(Ksiwx4 | Zn6wx4));
assign Wriwx4 = (Rsiwx4 & Ysiwx4);
assign Ysiwx4 = (Fdsvx4 | R89vx4);
assign Rsiwx4 = (K79vx4 | Fb9vx4);
assign Epiwx4 = (~(Ftiwx4 & Mtiwx4));
assign Mtiwx4 = (~(Q4wvx4 & Sjwvx4));
assign Ftiwx4 = (H5fwx4 | Qsewx4);
assign Bkiwx4 = (Ttiwx4 & Auiwx4);
assign Auiwx4 = (~(Huiwx4 & Efgvx4));
assign Ttiwx4 = (Ujxvx4 ? Vuiwx4 : Ouiwx4);
assign Vuiwx4 = (~(Cviwx4 & O76wx4));
assign Cviwx4 = (~(H33wx4 | E78wx4));
assign Ouiwx4 = (~(Jviwx4 & Qviwx4));
assign Qviwx4 = (!Qhqvx4);
assign Jviwx4 = (~(Xviwx4 | U0ovx4));
assign Fvhvx4 = (Ewiwx4 & Lwiwx4);
assign Lwiwx4 = (~(Swiwx4 & Zwiwx4));
assign Zwiwx4 = (Gxiwx4 & Nxiwx4);
assign Nxiwx4 = (Uxiwx4 & Byiwx4);
assign Byiwx4 = (Iyiwx4 & Pyiwx4);
assign Pyiwx4 = (~(Qsewx4 & Wyiwx4));
assign Wyiwx4 = (~(Dziwx4 & Kziwx4));
assign Kziwx4 = (~(Wvewx4 & Rziwx4));
assign Rziwx4 = (~(Yziwx4 & F0jwx4));
assign F0jwx4 = (M0jwx4 & Fdsvx4);
assign M0jwx4 = (W49vx4 | K79vx4);
assign Yziwx4 = (~(Y5svx4 | C1svx4));
assign Iyiwx4 = (~(Ahwvx4 & T0jwx4));
assign T0jwx4 = (~(A1jwx4 & H1jwx4));
assign H1jwx4 = (~(O1jwx4 & V1jwx4));
assign V1jwx4 = (~(C2jwx4 & J2jwx4));
assign J2jwx4 = (Qfsvx4 | K79vx4);
assign C2jwx4 = (~(Zn6wx4 | Y99vx4));
assign A1jwx4 = (Epxvx4 | Dj6wx4);
assign Uxiwx4 = (Q2jwx4 & X2jwx4);
assign X2jwx4 = (~(Z7fwx4 & E3jwx4));
assign E3jwx4 = (~(L3jwx4 & S3jwx4));
assign S3jwx4 = (~(Z3jwx4 & G4jwx4));
assign G4jwx4 = (N4jwx4 & Ujxvx4);
assign N4jwx4 = (Eiqvx4 | Auqvx4);
assign Auqvx4 = (~(W5yvx4 | Mcgvx4));
assign L3jwx4 = (O58wx4 | Msyvx4);
assign Q2jwx4 = (~(Fjewx4 & U4jwx4));
assign U4jwx4 = (~(B5jwx4 & I5jwx4));
assign I5jwx4 = (~(P5jwx4 & Qp3wx4));
assign B5jwx4 = (Jf6wx4 | B4dwx4);
assign Jf6wx4 = (!Nuewx4);
assign Gxiwx4 = (W5jwx4 & D6jwx4);
assign D6jwx4 = (K6jwx4 & R6jwx4);
assign R6jwx4 = (~(Y6jwx4 & Izwvx4));
assign Y6jwx4 = (~(F7jwx4 & Y2ovx4));
assign Y2ovx4 = (~(Ri7wx4 & U0ovx4));
assign F7jwx4 = (~(Jp3wx4 & Eznvx4));
assign K6jwx4 = (Pdqvx4 | Efgvx4);
assign Pdqvx4 = (!M7jwx4);
assign W5jwx4 = (T7jwx4 & A8jwx4);
assign A8jwx4 = (Kvfwx4 | Fjgvx4);
assign T7jwx4 = (H8jwx4 | Zg6wx4);
assign Zg6wx4 = (~(Ki8vx4 | Mj8vx4));
assign Swiwx4 = (O8jwx4 & V8jwx4);
assign V8jwx4 = (C9jwx4 & J9jwx4);
assign J9jwx4 = (Q9jwx4 & X9jwx4);
assign X9jwx4 = (Xhiwx4 | Mj8vx4);
assign Q9jwx4 = (~(Pcyvx4 & Eajwx4));
assign Eajwx4 = (~(Lajwx4 & Sajwx4));
assign Sajwx4 = (Y47wx4 | Wt2wx4);
assign Lajwx4 = (Zajwx4 & Gbjwx4);
assign Gbjwx4 = (Fscwx4 | Z6gvx4);
assign Zajwx4 = (Zj3wx4 | Bl3wx4);
assign C9jwx4 = (Nbjwx4 & Ubjwx4);
assign Ubjwx4 = (~(Sh9vx4 & Bcjwx4));
assign Bcjwx4 = (~(Icjwx4 & Pcjwx4));
assign Pcjwx4 = (Ct6wx4 | Icyvx4);
assign Icjwx4 = (Wcjwx4 & Ddjwx4);
assign Ddjwx4 = (~(Kdjwx4 & Jjgwx4));
assign Kdjwx4 = (~(Izwvx4 | Y99vx4));
assign Wcjwx4 = (~(U1fwx4 & Wvewx4));
assign Nbjwx4 = (~(A0zvx4 & Rdjwx4));
assign Rdjwx4 = (Ydjwx4 | Fejwx4);
assign Fejwx4 = (Bl3wx4 ? Hw2wx4 : B1ovx4);
assign Ydjwx4 = (Mejwx4 | U6hwx4);
assign U6hwx4 = (~(Msyvx4 | Dbgvx4));
assign Mejwx4 = (~(S87wx4 | Emewx4));
assign O8jwx4 = (Tejwx4 & Afjwx4);
assign Afjwx4 = (Hfjwx4 & Ofjwx4);
assign Ofjwx4 = (~(Vfjwx4 & Lcpvx4));
assign Vfjwx4 = (~(Cgjwx4 & Jgjwx4));
assign Jgjwx4 = (Qgjwx4 & Xgjwx4);
assign Xgjwx4 = (~(Soyvx4 & Qfsvx4));
assign Soyvx4 = (~(Izwvx4 | Sh9vx4));
assign Qgjwx4 = (Ehjwx4 & Lhjwx4);
assign Lhjwx4 = (~(Shjwx4 & O1jwx4));
assign Shjwx4 = (~(Izwvx4 | Dj6wx4));
assign Ehjwx4 = (~(Nkpvx4 & Zhjwx4));
assign Zhjwx4 = (Gijwx4 | Nijwx4);
assign Nijwx4 = (Uasvx4 ? Zn6wx4 : N3svx4);
assign Gijwx4 = (Uijwx4 | Txewx4);
assign Cgjwx4 = (Bjjwx4 & Ijjwx4);
assign Ijjwx4 = (X5gwx4 | Fdsvx4);
assign Bjjwx4 = (Yj6wx4 | Sh9vx4);
assign Hfjwx4 = (~(Howvx4 & Nv6wx4));
assign Tejwx4 = (~(Pjjwx4 | Q6fwx4));
assign Q6fwx4 = (~(Wjjwx4 & Dkjwx4));
assign Dkjwx4 = (Kkjwx4 & Svyvx4);
assign Kkjwx4 = (~(Ccovx4 | Oowvx4));
assign Oowvx4 = (~(M1xvx4 | Izwvx4));
assign Wjjwx4 = (Rkjwx4 & Ykjwx4);
assign Ykjwx4 = (~(Fljwx4 & Dmgvx4));
assign Fljwx4 = (~(S4xvx4 | Efgvx4));
assign Pjjwx4 = (Qfsvx4 ? Pswvx4 : Mljwx4);
assign Ewiwx4 = (U9gvx4 | hready_i);
assign Yuhvx4 = (!Tljwx4);
assign Tljwx4 = (Ccovx4 ? F3ovx4 : Amjwx4);
assign Amjwx4 = (Hmjwx4 & Omjwx4);
assign Omjwx4 = (Vmjwx4 & Cnjwx4);
assign Cnjwx4 = (Jnjwx4 & Qnjwx4);
assign Qnjwx4 = (Xnjwx4 & Sygwx4);
assign Sygwx4 = (~(Eojwx4 & Srgwx4));
assign Eojwx4 = (~(Bl3wx4 | Z6gvx4));
assign Jnjwx4 = (Svyvx4 & Og4wx4);
assign Vmjwx4 = (Lojwx4 & Sojwx4);
assign Sojwx4 = (~(Zojwx4 & Q5gvx4));
assign Zojwx4 = (~(Sznvx4 | K7xvx4));
assign Lojwx4 = (Gpjwx4 & Fhgwx4);
assign Gpjwx4 = (~(Npjwx4 & Gh6wx4));
assign Npjwx4 = (~(Zjwvx4 | Bzwvx4));
assign Bzwvx4 = (~(Qfsvx4 | Xmsvx4));
assign Hmjwx4 = (Upjwx4 & Bqjwx4);
assign Bqjwx4 = (Iqjwx4 & Pqjwx4);
assign Pqjwx4 = (Qhqvx4 | Wqjwx4);
assign Iqjwx4 = (Drjwx4 & Krjwx4);
assign Krjwx4 = (~(Rrjwx4 & M3ovx4));
assign Rrjwx4 = (~(Yrjwx4 & Fsjwx4));
assign Fsjwx4 = (F57wx4 | Zrvvx4);
assign Yrjwx4 = (Msjwx4 & Tsjwx4);
assign Tsjwx4 = (~(Atjwx4 & P9fwx4));
assign Atjwx4 = (~(O4ovx4 | Vdgvx4));
assign Msjwx4 = (Efewx4 | A8yvx4);
assign Drjwx4 = (~(Htjwx4 & R7qvx4));
assign Htjwx4 = (~(Otjwx4 & Vtjwx4));
assign Vtjwx4 = (Cujwx4 & Jujwx4);
assign Jujwx4 = (Qujwx4 & Xujwx4);
assign Xujwx4 = (~(Evjwx4 & V1yvx4));
assign Evjwx4 = (Lvjwx4 & M1xvx4);
assign Lvjwx4 = (~(Svjwx4 & Zvjwx4));
assign Zvjwx4 = (~(Gwjwx4 & Qfsvx4));
assign Gwjwx4 = (~(Nwjwx4 & R3fwx4));
assign R3fwx4 = (Uwjwx4 & Bxjwx4);
assign Bxjwx4 = (~(Ixjwx4 & Fb9vx4));
assign Ixjwx4 = (~(Y5svx4 | Y99vx4));
assign Uwjwx4 = (~(Mc9vx4 & Pxjwx4));
assign Pxjwx4 = (Y99vx4 | Ugewx4);
assign Nwjwx4 = (Sh9vx4 & Wxjwx4);
assign Wxjwx4 = (Tc7wx4 | J16wx4);
assign Tc7wx4 = (!Ix5wx4);
assign Svjwx4 = (~(Txewx4 & Hh3wx4));
assign Qujwx4 = (~(Dyjwx4 & Kg9vx4));
assign Dyjwx4 = (Ud9vx4 & Kyjwx4);
assign Kyjwx4 = (~(Ryjwx4 & Yyjwx4));
assign Yyjwx4 = (~(Fzjwx4 & Mzjwx4));
assign Mzjwx4 = (Tzjwx4 & Wvewx4);
assign Tzjwx4 = (~(D69vx4 | K79vx4));
assign Fzjwx4 = (A0kwx4 & Qxgwx4);
assign A0kwx4 = (O1jwx4 & Hyewx4);
assign Ryjwx4 = (Ulgwx4 | H0kwx4);
assign Cujwx4 = (O0kwx4 & V0kwx4);
assign V0kwx4 = (~(C1kwx4 & O1jwx4));
assign C1kwx4 = (~(Ct6wx4 | H5fwx4));
assign O0kwx4 = (~(J1kwx4 & Howvx4));
assign J1kwx4 = (~(Mv2wx4 | U9gvx4));
assign Otjwx4 = (Q1kwx4 & X1kwx4);
assign X1kwx4 = (E2kwx4 & L2kwx4);
assign L2kwx4 = (~(Wnfwx4 & A0zvx4));
assign Wnfwx4 = (~(S87wx4 | Fjewx4));
assign E2kwx4 = (~(Sjwvx4 & S2kwx4));
assign S2kwx4 = (~(Z2kwx4 & G3kwx4));
assign Z2kwx4 = (N3kwx4 & U3kwx4);
assign U3kwx4 = (~(B4kwx4 & Pyxvx4));
assign B4kwx4 = (Ud9vx4 ? Dj6wx4 : Uasvx4);
assign N3kwx4 = (X5gwx4 | Abgwx4);
assign Q1kwx4 = (I4kwx4 & P4kwx4);
assign P4kwx4 = (~(Oigwx4 & Wshwx4));
assign I4kwx4 = (Keqvx4 | K7xvx4);
assign Upjwx4 = (W4kwx4 & D5kwx4);
assign D5kwx4 = (Us2wx4 ? R5kwx4 : K5kwx4);
assign R5kwx4 = (Gjxvx4 | Nggvx4);
assign K5kwx4 = (~(Vdgvx4 & Y5kwx4));
assign Y5kwx4 = (~(Pxyvx4 & Lg6wx4));
assign Lg6wx4 = (~(Mj8vx4 & Kzxvx4));
assign W4kwx4 = (H2xvx4 & F6kwx4);
assign F6kwx4 = (Njxvx4 | Whgvx4);
assign Ruhvx4 = (M6kwx4 & T6kwx4);
assign T6kwx4 = (~(A7kwx4 & H7kwx4));
assign H7kwx4 = (O7kwx4 & V7kwx4);
assign V7kwx4 = (C8kwx4 & J8kwx4);
assign J8kwx4 = (Q8kwx4 & X8kwx4);
assign Q8kwx4 = (~(E9kwx4 & Os6wx4));
assign Os6wx4 = (~(D69vx4 | R89vx4));
assign E9kwx4 = (~(Bhewx4 | L9kwx4));
assign L9kwx4 = (~(Ryrvx4 | N3svx4));
assign Bhewx4 = (~(S9kwx4 & Z9kwx4));
assign Z9kwx4 = (~(Gakwx4 | J8svx4));
assign Gakwx4 = (!Blwvx4);
assign Blwvx4 = (~(Abgwx4 | Qfsvx4));
assign S9kwx4 = (Hyewx4 & N9ewx4);
assign Hyewx4 = (Nakwx4 & Uakwx4);
assign Uakwx4 = (~(I29vx4 | P39vx4));
assign C8kwx4 = (Bbkwx4 & Ibkwx4);
assign Ibkwx4 = (~(Pbkwx4 & Wbkwx4));
assign Pbkwx4 = (Keiwx4 & Howvx4);
assign Bbkwx4 = (~(Dckwx4 & Lxwvx4));
assign Dckwx4 = (Qaqvx4 & Kckwx4);
assign Kckwx4 = (~(Rckwx4 & Yckwx4));
assign Yckwx4 = (~(Fdkwx4 & O3hwx4));
assign Fdkwx4 = (~(Uasvx4 | Dfpvx4));
assign Rckwx4 = (Xmsvx4 | Bisvx4);
assign O7kwx4 = (Mdkwx4 & Tdkwx4);
assign Tdkwx4 = (Aekwx4 & Hekwx4);
assign Hekwx4 = (~(Oekwx4 & Gh6wx4));
assign Oekwx4 = (Vekwx4 & O4ovx4);
assign Vekwx4 = (~(G3kwx4 & Cfkwx4));
assign Cfkwx4 = (~(Jfkwx4 & Ahwvx4));
assign Jfkwx4 = (Hh3wx4 & J8svx4);
assign Hh3wx4 = (Fdsvx4 & Qfsvx4);
assign G3kwx4 = (Dziwx4 | Dfpvx4);
assign Aekwx4 = (~(Qfkwx4 & Xfkwx4));
assign Qfkwx4 = (~(K7xvx4 | Vdgvx4));
assign Mdkwx4 = (Egkwx4 & Lgkwx4);
assign Lgkwx4 = (~(Sgkwx4 & Mcewx4));
assign Sgkwx4 = (~(Oedwx4 | F3ovx4));
assign Egkwx4 = (~(Z9dwx4 & Zgkwx4));
assign Zgkwx4 = (Liqvx4 | Mcewx4);
assign A7kwx4 = (Ghkwx4 & Nhkwx4);
assign Nhkwx4 = (Uhkwx4 & Bikwx4);
assign Bikwx4 = (Iikwx4 & Pikwx4);
assign Pikwx4 = (~(Wdxvx4 & Wikwx4));
assign Wikwx4 = (~(Djkwx4 & Kjkwx4));
assign Kjkwx4 = (Gjxvx4 | S4xvx4);
assign Djkwx4 = (~(O76wx4 & Efgvx4));
assign Iikwx4 = (~(Su6wx4 & C2yvx4));
assign Su6wx4 = (Rjkwx4 & Yjkwx4);
assign Yjkwx4 = (K8hwx4 & Bl3wx4);
assign Rjkwx4 = (W7hwx4 & Cjgwx4);
assign Cjgwx4 = (Howvx4 & Kngwx4);
assign Uhkwx4 = (Fkkwx4 & Mkkwx4);
assign Mkkwx4 = (~(Fjewx4 & Tkkwx4));
assign Tkkwx4 = (~(Alkwx4 & Hlkwx4));
assign Hlkwx4 = (~(Gs2wx4 & Qp3wx4));
assign Gs2wx4 = (Jp3wx4 & O4ovx4);
assign Alkwx4 = (Olkwx4 & Vlkwx4);
assign Vlkwx4 = (~(Cmkwx4 & Jmkwx4));
assign Jmkwx4 = (~(Jppvx4 | Z6gvx4));
assign Cmkwx4 = (~(Qmkwx4 | Xp3wx4));
assign Xp3wx4 = (!U63wx4);
assign U63wx4 = (~(Oedwx4 | Mcgvx4));
assign Olkwx4 = (~(O76wx4 & Xmkwx4));
assign Xmkwx4 = (~(Chxvx4 & Enkwx4));
assign Enkwx4 = (Gcqvx4 | U9gvx4);
assign Chxvx4 = (Hq1wx4 | Us2wx4);
assign Fkkwx4 = (~(Lnkwx4 & R7qvx4));
assign Lnkwx4 = (~(Snkwx4 & Znkwx4));
assign Znkwx4 = (Gokwx4 & Ej3wx4);
assign Ej3wx4 = (~(Nokwx4 & Ukpvx4));
assign Nokwx4 = (Pswvx4 & Abgwx4);
assign Gokwx4 = (~(Uokwx4 & Bpkwx4));
assign Bpkwx4 = (~(Ud9vx4 | Sh9vx4));
assign Uokwx4 = (~(Xaxvx4 | Ho8vx4));
assign Xaxvx4 = (!Ipkwx4);
assign Snkwx4 = (Ppkwx4 & Wpkwx4);
assign Wpkwx4 = (~(Dqkwx4 & Ukpvx4));
assign Dqkwx4 = (~(Oohwx4 | J8svx4));
assign Oohwx4 = (!Pswvx4);
assign Ppkwx4 = (Pxyvx4 | S4xvx4);
assign Ghkwx4 = (Kqkwx4 & Rqkwx4);
assign Rqkwx4 = (Uv6wx4 & V76wx4);
assign V76wx4 = (Yqkwx4 & Frkwx4);
assign Frkwx4 = (Zq3wx4 | Nggvx4);
assign Zq3wx4 = (~(A0zvx4 & B73wx4));
assign Yqkwx4 = (Mrkwx4 & Gwyvx4);
assign Gwyvx4 = (O58wx4 | Gjxvx4);
assign O58wx4 = (!Ptgwx4);
assign Uv6wx4 = (Trkwx4 & Fhgwx4);
assign Trkwx4 = (~(Ccovx4 | M7jwx4));
assign M7jwx4 = (~(A8yvx4 | S4xvx4));
assign A8yvx4 = (!Zzfwx4);
assign Kqkwx4 = (Askwx4 & Unewx4);
assign Unewx4 = (Hskwx4 & Oskwx4);
assign Oskwx4 = (~(V06wx4 & J16wx4));
assign V06wx4 = (N9ewx4 & A4gwx4);
assign Hskwx4 = (Vskwx4 & Ctkwx4);
assign Ctkwx4 = (~(Jtkwx4 & Mcewx4));
assign Mcewx4 = (B73wx4 & Pcyvx4);
assign Vskwx4 = (~(N9ewx4 & Bisvx4));
assign N9ewx4 = (Gh6wx4 & Ohwvx4);
assign Gh6wx4 = (Aj9vx4 & R7qvx4);
assign Askwx4 = (Xmsvx4 ? Xtkwx4 : Qtkwx4);
assign Xtkwx4 = (~(Eukwx4 & X16wx4));
assign Eukwx4 = (Ud9vx4 & Lukwx4);
assign Lukwx4 = (~(Zjwvx4 & Sukwx4));
assign Sukwx4 = (~(Ix5wx4 & Xhxvx4));
assign Qtkwx4 = (~(Px5wx4 & Zukwx4));
assign Zukwx4 = (~(Gvkwx4 & Nvkwx4));
assign Nvkwx4 = (~(Qxgwx4 | Ix5wx4));
assign Ix5wx4 = (~(Mc9vx4 | Fb9vx4));
assign Qxgwx4 = (Uvkwx4 & G27wx4);
assign Uvkwx4 = (~(J8svx4 | R89vx4));
assign Gvkwx4 = (Bwkwx4 & Iwkwx4);
assign Iwkwx4 = (~(Pwkwx4 & R89vx4));
assign Pwkwx4 = (~(Txewx4 | Mc9vx4));
assign Txewx4 = (~(K79vx4 | Y99vx4));
assign Bwkwx4 = (~(Ugewx4 & Tr6wx4));
assign Ugewx4 = (Wwkwx4 & Lwxvx4);
assign Lwxvx4 = (Uz8vx4 & B19vx4);
assign Wwkwx4 = (~(Vtrvx4 | Y5svx4));
assign Vtrvx4 = (!I29vx4);
assign Px5wx4 = (Dxkwx4 & X16wx4);
assign X16wx4 = (Mgwvx4 & Qaqvx4);
assign Dxkwx4 = (~(Dziwx4 | Kg9vx4));
assign M6kwx4 = (Vdgvx4 | hready_i);
assign Kuhvx4 = (K6yvx4 ? Kxkwx4 : Xq8vx4);
assign Kxkwx4 = (~(Rxkwx4 & Yxkwx4));
assign Yxkwx4 = (Fykwx4 & Mykwx4);
assign Mykwx4 = (~(P39vx4 & Zayvx4));
assign Fykwx4 = (Tykwx4 & Azkwx4);
assign Azkwx4 = (~(H8yvx4 & Uz8vx4));
assign Tykwx4 = (~(C9yvx4 & Hzkwx4));
assign Hzkwx4 = (~(Ozkwx4 & Vzkwx4));
assign Vzkwx4 = (C0lwx4 & J0lwx4);
assign J0lwx4 = (Q0lwx4 | Emewx4);
assign C0lwx4 = (~(X0lwx4 & X9yvx4));
assign Ozkwx4 = (E1lwx4 & L1lwx4);
assign L1lwx4 = (~(Sayvx4 & S1lwx4));
assign E1lwx4 = (~(Su9vx4 & G6wvx4));
assign Rxkwx4 = (Z1lwx4 & G2lwx4);
assign Z1lwx4 = (N2lwx4 & U2lwx4);
assign U2lwx4 = (Icyvx4 | N3svx4);
assign N2lwx4 = (~(Ot9vx4 & Pcyvx4));
assign Duhvx4 = (~(B3lwx4 & I3lwx4));
assign I3lwx4 = (P3lwx4 & W3lwx4);
assign W3lwx4 = (~(Xdfwx4 & Dmh2z4[24]));
assign P3lwx4 = (D4lwx4 & Lefwx4);
assign D4lwx4 = (Sefwx4 | O3pvx4);
assign O3pvx4 = (K4lwx4 & R4lwx4);
assign R4lwx4 = (Y4lwx4 & F5lwx4);
assign F5lwx4 = (~(W6iwx4 & Hmyvx4));
assign Y4lwx4 = (M5lwx4 & R7iwx4);
assign M5lwx4 = (~(Pjyvx4 & F8iwx4));
assign K4lwx4 = (T5lwx4 & A6lwx4);
assign A6lwx4 = (~(Rkyvx4 & H9iwx4));
assign T5lwx4 = (~(Tlyvx4 & V9iwx4));
assign B3lwx4 = (H6lwx4 & O6lwx4);
assign O6lwx4 = (~(Roh2z4[23] & Mifwx4));
assign H6lwx4 = (~(vis_pc_o[23] & Qaiwx4));
assign Wthvx4 = (~(V6lwx4 & C7lwx4));
assign C7lwx4 = (J7lwx4 & Q7lwx4);
assign Q7lwx4 = (~(Xdfwx4 & Dmh2z4[31]));
assign J7lwx4 = (X7lwx4 & Lefwx4);
assign X7lwx4 = (Sefwx4 | R5zvx4);
assign R5zvx4 = (E8lwx4 & L8lwx4);
assign L8lwx4 = (S8lwx4 & Z8lwx4);
assign Z8lwx4 = (~(G9lwx4 & V9iwx4));
assign S8lwx4 = (N9lwx4 & R7iwx4);
assign N9lwx4 = (~(W6iwx4 & U9lwx4));
assign E8lwx4 = (Balwx4 & Ialwx4);
assign Ialwx4 = (~(Palwx4 & H9iwx4));
assign Balwx4 = (~(Walwx4 & F8iwx4));
assign V6lwx4 = (Dblwx4 & Kblwx4);
assign Kblwx4 = (~(Roh2z4[30] & Mifwx4));
assign Dblwx4 = (~(vis_pc_o[30] & Qaiwx4));
assign Pthvx4 = (Yafwx4 ? Rblwx4 : Tjh2z4[1]);
assign Rblwx4 = (~(Yblwx4 & Fclwx4));
assign Fclwx4 = (Mclwx4 & Tclwx4);
assign Tclwx4 = (~(Q3iwx4 & W49vx4));
assign Mclwx4 = (Adlwx4 & Hdlwx4);
assign Hdlwx4 = (~(Odlwx4 & Vdlwx4));
assign Vdlwx4 = (~(U4yvx4 | Ud9vx4));
assign Odlwx4 = (Kg9vx4 & K8hwx4);
assign Adlwx4 = (Uasvx4 | J3iwx4);
assign Yblwx4 = (Celwx4 & Jelwx4);
assign Jelwx4 = (~(B19vx4 & E4iwx4));
assign Ithvx4 = (~(Qelwx4 & Xelwx4));
assign Xelwx4 = (Eflwx4 & Lflwx4);
assign Lflwx4 = (~(Roh2z4[18] & Mifwx4));
assign Eflwx4 = (Sflwx4 & Zflwx4);
assign Zflwx4 = (Sefwx4 | Bo0wx4);
assign Bo0wx4 = (Gglwx4 & Nglwx4);
assign Nglwx4 = (Uglwx4 & Bhlwx4);
assign Bhlwx4 = (~(W6iwx4 & Ihlwx4));
assign Uglwx4 = (~(Phlwx4 & Whlwx4));
assign Gglwx4 = (Dilwx4 & Kilwx4);
assign Kilwx4 = (~(Rilwx4 & Yilwx4));
assign Dilwx4 = (~(Fjlwx4 & Mjlwx4));
assign Sflwx4 = (~(Xdfwx4 & Dmh2z4[19]));
assign Qelwx4 = (Tjlwx4 & Aklwx4);
assign Aklwx4 = (~(vis_pc_o[18] & Qaiwx4));
assign Bthvx4 = (~(Hklwx4 & Oklwx4));
assign Oklwx4 = (~(Vklwx4 & Cllwx4));
assign Hklwx4 = (Qllwx4 ? Jllwx4 : Xy8wx4);
assign Jllwx4 = (Xllwx4 & Emlwx4);
assign Emlwx4 = (Lmlwx4 & Smlwx4);
assign Smlwx4 = (Nrwvx4 & Bswvx4);
assign Nrwvx4 = (~(R5dwx4 & Fjgvx4));
assign Lmlwx4 = (Zmlwx4 & Gnlwx4);
assign Gnlwx4 = (~(Nnlwx4 & Mc9vx4));
assign Nnlwx4 = (Unlwx4 & Lcpvx4);
assign Unlwx4 = (~(O1yvx4 & Bolwx4));
assign Bolwx4 = (~(Xhxvx4 & C2yvx4));
assign O1yvx4 = (~(Uuewx4 & O4ovx4));
assign Uuewx4 = (Qsewx4 & Cn8vx4);
assign Zmlwx4 = (~(Iolwx4 & Polwx4));
assign Polwx4 = (Ceewx4 ^ Jeewx4);
assign Jeewx4 = (Anxvx4 | U5bwx4);
assign Anxvx4 = (~(H9xvx4 & Qm9vx4));
assign Ceewx4 = (~(Yo9vx4 & Zrvvx4));
assign Iolwx4 = (Vopvx4 & Jj9wx4);
assign Vopvx4 = (~(Wolwx4 & Dplwx4));
assign Wolwx4 = (Kplwx4 & Rplwx4);
assign Rplwx4 = (Yplwx4 | Us2wx4);
assign Kplwx4 = (~(Ilpvx4 & Fqlwx4));
assign Xllwx4 = (Mqlwx4 & Tqlwx4);
assign Tqlwx4 = (Arlwx4 & Hrlwx4);
assign Hrlwx4 = (~(Orlwx4 & Vsevx4));
assign Arlwx4 = (~(W49vx4 & Vrlwx4));
assign Mqlwx4 = (Cslwx4 & Jslwx4);
assign Jslwx4 = (~(Dsqvx4 & Fb9vx4));
assign Cslwx4 = (~(P39vx4 & Qslwx4));
assign Ushvx4 = (~(Xslwx4 & Etlwx4));
assign Etlwx4 = (~(Fjgvx4 & Ltlwx4));
assign Ltlwx4 = (~(Stlwx4 & Ztlwx4));
assign Ztlwx4 = (Dmgvx4 | Efgvx4);
assign Stlwx4 = (~(Ccovx4 | Ptgwx4));
assign Ptgwx4 = (~(Mcgvx4 | Whgvx4));
assign Xslwx4 = (~(Gulwx4 & hready_i));
assign Gulwx4 = (~(Nulwx4 & Uulwx4));
assign Uulwx4 = (Bvlwx4 & Ivlwx4);
assign Ivlwx4 = (~(Msyvx4 & Pvlwx4));
assign Pvlwx4 = (~(Wvlwx4 & Dwlwx4));
assign Dwlwx4 = (~(Kwlwx4 & Z7fwx4));
assign Kwlwx4 = (~(Dbgvx4 | Whgvx4));
assign Wvlwx4 = (Bqcwx4 | Tv2wx4);
assign Bqcwx4 = (!A0zvx4);
assign Bvlwx4 = (Rwlwx4 & Bswvx4);
assign Rwlwx4 = (~(Ywlwx4 & Ho8vx4));
assign Ywlwx4 = (Sh9vx4 & Fxlwx4);
assign Fxlwx4 = (~(Bdqvx4 & Mxlwx4));
assign Mxlwx4 = (~(Wbkwx4 & Y38wx4));
assign Y38wx4 = (~(S4xvx4 | Fjgvx4));
assign Nulwx4 = (Txlwx4 & Aylwx4);
assign Aylwx4 = (S87wx4 | O4ovx4);
assign Txlwx4 = (U36wx4 & Hylwx4);
assign Hylwx4 = (Sznvx4 | Z9dwx4);
assign U36wx4 = (Gjxvx4 | Hq1wx4);
assign Nshvx4 = (J5vvx4 ? By4wx4 : Q5gvx4);
assign By4wx4 = (Xlevx4 & Oylwx4);
assign Oylwx4 = (~(Vylwx4 & Czlwx4));
assign Czlwx4 = (Jzlwx4 & Qzlwx4);
assign Qzlwx4 = (~(Jyevx4 | Tzevx4));
assign Jzlwx4 = (~(Pvevx4 | Zwevx4));
assign Vylwx4 = (Xzlwx4 & E0mwx4);
assign E0mwx4 = (~(Z3fvx4 | K5fvx4));
assign Xzlwx4 = (~(D1fvx4 | O2fvx4));
assign Gshvx4 = (hready_i ? hwrite_o : Pp8vx4);
assign hwrite_o = (~(L0mwx4 & S0mwx4));
assign S0mwx4 = (Z0mwx4 & G1mwx4);
assign G1mwx4 = (~(Pa7wx4 & N1mwx4));
assign N1mwx4 = (~(Qhqvx4 & U1mwx4));
assign U1mwx4 = (~(B2mwx4 & Ucqvx4));
assign B2mwx4 = (B73wx4 & R7qvx4);
assign Qhqvx4 = (~(Kzxvx4 & S4xvx4));
assign L0mwx4 = (I2mwx4 & P2mwx4);
assign P2mwx4 = (~(B1vvx4 & W2mwx4));
assign W2mwx4 = (~(Jrnvx4 & D3mwx4));
assign D3mwx4 = (~(K3mwx4 & Fqlwx4));
assign K3mwx4 = (~(Oedwx4 | Mvgwx4));
assign Jrnvx4 = (!Vhpvx4);
assign Vhpvx4 = (~(Oedwx4 | Zrvvx4));
assign Zrhvx4 = (hready_i ? R3mwx4 : Hx8vx4);
assign R3mwx4 = (~(Y3mwx4 & F4mwx4));
assign F4mwx4 = (~(M4mwx4 & T4mwx4));
assign T4mwx4 = (Pcyvx4 & X43wx4);
assign M4mwx4 = (~(Mvgwx4 | Mv2wx4));
assign Y3mwx4 = (~(A5mwx4 & H5mwx4));
assign A5mwx4 = (B73wx4 & Vdgvx4);
assign Srhvx4 = (J5vvx4 ? Ye4wx4 : Rkgvx4);
assign J5vvx4 = (Fjgvx4 & hready_i);
assign Lrhvx4 = (!O5mwx4);
assign O5mwx4 = (Ccovx4 ? Efewx4 : V5mwx4);
assign V5mwx4 = (~(C6mwx4 | J6mwx4));
assign J6mwx4 = (~(Q6mwx4 | F3vvx4));
assign Erhvx4 = (!X6mwx4);
assign X6mwx4 = (hready_i ? E7mwx4 : Neovx4);
assign Xqhvx4 = (Bpsvx4 ? Xcovx4 : Mxfvx4);
assign Xcovx4 = (!Ueovx4);
assign Qqhvx4 = (~(L7mwx4 & S7mwx4));
assign S7mwx4 = (~(Z7mwx4 & hrdata_i[16]));
assign L7mwx4 = (~(Cbfvx4 & Sorvx4));
assign Jqhvx4 = (~(G8mwx4 & N8mwx4));
assign N8mwx4 = (~(Z7mwx4 & hrdata_i[17]));
assign G8mwx4 = (~(Mcfvx4 & Sorvx4));
assign Cqhvx4 = (~(U8mwx4 & B9mwx4));
assign B9mwx4 = (~(Z7mwx4 & hrdata_i[18]));
assign U8mwx4 = (~(Wdfvx4 & Sorvx4));
assign Vphvx4 = (~(I9mwx4 & P9mwx4));
assign P9mwx4 = (~(Z7mwx4 & hrdata_i[19]));
assign I9mwx4 = (~(Gffvx4 & Sorvx4));
assign Ophvx4 = (~(W9mwx4 & Damwx4));
assign Damwx4 = (~(Z7mwx4 & hrdata_i[20]));
assign W9mwx4 = (~(Qgfvx4 & Sorvx4));
assign Hphvx4 = (~(Kamwx4 & Ramwx4));
assign Ramwx4 = (~(Z7mwx4 & hrdata_i[21]));
assign Kamwx4 = (~(Aifvx4 & Sorvx4));
assign Aphvx4 = (~(Yamwx4 & Fbmwx4));
assign Fbmwx4 = (~(Z7mwx4 & hrdata_i[22]));
assign Yamwx4 = (~(Kjfvx4 & Sorvx4));
assign Tohvx4 = (~(Mbmwx4 & Tbmwx4));
assign Tbmwx4 = (~(Z7mwx4 & hrdata_i[23]));
assign Mbmwx4 = (~(Ukfvx4 & Sorvx4));
assign Mohvx4 = (~(Acmwx4 & Hcmwx4));
assign Hcmwx4 = (~(Z7mwx4 & hrdata_i[24]));
assign Acmwx4 = (~(Emfvx4 & Sorvx4));
assign Fohvx4 = (~(Ocmwx4 & Vcmwx4));
assign Vcmwx4 = (~(Z7mwx4 & hrdata_i[25]));
assign Ocmwx4 = (~(Onfvx4 & Sorvx4));
assign Ynhvx4 = (~(Cdmwx4 & Jdmwx4));
assign Jdmwx4 = (~(Z7mwx4 & hrdata_i[26]));
assign Cdmwx4 = (~(Yofvx4 & Sorvx4));
assign Rnhvx4 = (~(Qdmwx4 & Xdmwx4));
assign Xdmwx4 = (~(Z7mwx4 & hrdata_i[27]));
assign Qdmwx4 = (~(Jqfvx4 & Sorvx4));
assign Knhvx4 = (~(Eemwx4 & Lemwx4));
assign Lemwx4 = (~(Z7mwx4 & hrdata_i[28]));
assign Eemwx4 = (~(Urfvx4 & Sorvx4));
assign Dnhvx4 = (~(Semwx4 & Zemwx4));
assign Zemwx4 = (~(Z7mwx4 & hrdata_i[29]));
assign Semwx4 = (~(Ftfvx4 & Sorvx4));
assign Wmhvx4 = (~(Gfmwx4 & Nfmwx4));
assign Nfmwx4 = (~(Z7mwx4 & hrdata_i[30]));
assign Gfmwx4 = (~(Qufvx4 & Sorvx4));
assign Pmhvx4 = (~(Ufmwx4 & Bgmwx4));
assign Bgmwx4 = (~(Z7mwx4 & hrdata_i[31]));
assign Z7mwx4 = (Ueovx4 & Bpsvx4);
assign Ueovx4 = (Igmwx4 & vis_tbit_o);
assign Igmwx4 = (~(hresp_i | H0gvx4));
assign Ufmwx4 = (~(Bwfvx4 & Sorvx4));
assign Sorvx4 = (!Bpsvx4);
assign Bpsvx4 = (~(Neovx4 | Ccovx4));
assign Neovx4 = (!Xyfvx4);
assign Imhvx4 = (~(Pgmwx4 & Wgmwx4));
assign Wgmwx4 = (Dhmwx4 & Khmwx4);
assign Khmwx4 = (~(Xdfwx4 & Dmh2z4[2]));
assign Dhmwx4 = (Rhmwx4 & Lefwx4);
assign Rhmwx4 = (Sefwx4 | Zluvx4);
assign Zluvx4 = (Yhmwx4 & Fimwx4);
assign Fimwx4 = (Mimwx4 & Timwx4);
assign Timwx4 = (~(Ajmwx4 & Wjyvx4));
assign Mimwx4 = (Hjmwx4 & Kkyvx4);
assign Hjmwx4 = (~(Ojmwx4 & Amyvx4));
assign Yhmwx4 = (Vjmwx4 & Ckmwx4);
assign Ckmwx4 = (~(Jkmwx4 & Ykyvx4));
assign Vjmwx4 = (~(Qkmwx4 & Omyvx4));
assign Pgmwx4 = (Xkmwx4 & Elmwx4);
assign Elmwx4 = (~(Roh2z4[1] & Mifwx4));
assign Xkmwx4 = (Pnnvx4 | G6pvx4);
assign Pnnvx4 = (!vis_pc_o[1]);
assign Bmhvx4 = (~(Llmwx4 & Slmwx4));
assign Slmwx4 = (Zlmwx4 & Gmmwx4);
assign Gmmwx4 = (~(Xdfwx4 & Dmh2z4[3]));
assign Zlmwx4 = (Nmmwx4 & Lefwx4);
assign Nmmwx4 = (Sefwx4 | U0vvx4);
assign U0vvx4 = (Ummwx4 & Bnmwx4);
assign Bnmwx4 = (Inmwx4 & Pnmwx4);
assign Pnmwx4 = (~(Rilwx4 & Wjyvx4));
assign Inmwx4 = (Wnmwx4 & Kkyvx4);
assign Wnmwx4 = (~(Mjlwx4 & Ykyvx4));
assign Ummwx4 = (Domwx4 & Komwx4);
assign Komwx4 = (~(Whlwx4 & Omyvx4));
assign Domwx4 = (~(Ihlwx4 & Amyvx4));
assign Llmwx4 = (Romwx4 & Yomwx4);
assign Yomwx4 = (~(Roh2z4[2] & Mifwx4));
assign Romwx4 = (Fpmwx4 | G6pvx4);
assign Ulhvx4 = (~(Mpmwx4 & Tpmwx4));
assign Tpmwx4 = (Aqmwx4 & Hqmwx4);
assign Hqmwx4 = (~(Xdfwx4 & Dmh2z4[4]));
assign Aqmwx4 = (Oqmwx4 & Lefwx4);
assign Oqmwx4 = (Sefwx4 | Leuvx4);
assign Leuvx4 = (Vqmwx4 & Crmwx4);
assign Crmwx4 = (Jrmwx4 & Qrmwx4);
assign Qrmwx4 = (~(Xrmwx4 & Omyvx4));
assign Jrmwx4 = (Esmwx4 & Kkyvx4);
assign Esmwx4 = (~(Lsmwx4 & Ykyvx4));
assign Vqmwx4 = (Ssmwx4 & Zsmwx4);
assign Zsmwx4 = (~(Gtmwx4 & Amyvx4));
assign Ssmwx4 = (~(Ntmwx4 & Wjyvx4));
assign Mpmwx4 = (Utmwx4 & Bumwx4);
assign Bumwx4 = (~(Roh2z4[3] & Mifwx4));
assign Utmwx4 = (~(vis_pc_o[3] & Qaiwx4));
assign Nlhvx4 = (~(Iumwx4 & Pumwx4));
assign Pumwx4 = (Wumwx4 & Dvmwx4);
assign Dvmwx4 = (~(Xdfwx4 & Dmh2z4[5]));
assign Wumwx4 = (Kvmwx4 & Lefwx4);
assign Kvmwx4 = (Sefwx4 | Vcuvx4);
assign Vcuvx4 = (Rvmwx4 & Yvmwx4);
assign Yvmwx4 = (Fwmwx4 & Mwmwx4);
assign Mwmwx4 = (~(Twmwx4 & Omyvx4));
assign Fwmwx4 = (Axmwx4 & Kkyvx4);
assign Axmwx4 = (~(Hxmwx4 & Ykyvx4));
assign Rvmwx4 = (Oxmwx4 & Vxmwx4);
assign Vxmwx4 = (~(Cymwx4 & Amyvx4));
assign Oxmwx4 = (~(Jymwx4 & Wjyvx4));
assign Iumwx4 = (Qymwx4 & Xymwx4);
assign Xymwx4 = (~(Roh2z4[4] & Mifwx4));
assign Qymwx4 = (~(vis_pc_o[4] & Qaiwx4));
assign Glhvx4 = (~(Ezmwx4 & Lzmwx4));
assign Lzmwx4 = (Szmwx4 & Zzmwx4);
assign Zzmwx4 = (~(Xdfwx4 & Dmh2z4[6]));
assign Szmwx4 = (G0nwx4 & Lefwx4);
assign G0nwx4 = (Sefwx4 | Zuzvx4);
assign Zuzvx4 = (N0nwx4 & U0nwx4);
assign U0nwx4 = (B1nwx4 & I1nwx4);
assign I1nwx4 = (~(Y7iwx4 & Wjyvx4));
assign B1nwx4 = (P1nwx4 & Kkyvx4);
assign P1nwx4 = (~(O9iwx4 & Amyvx4));
assign N0nwx4 = (W1nwx4 & D2nwx4);
assign D2nwx4 = (~(A9iwx4 & Ykyvx4));
assign W1nwx4 = (~(D7iwx4 & Omyvx4));
assign Ezmwx4 = (K2nwx4 & R2nwx4);
assign R2nwx4 = (~(Roh2z4[5] & Mifwx4));
assign K2nwx4 = (~(vis_pc_o[5] & Qaiwx4));
assign Zkhvx4 = (~(Y2nwx4 & F3nwx4));
assign F3nwx4 = (M3nwx4 & T3nwx4);
assign T3nwx4 = (~(Xdfwx4 & Dmh2z4[7]));
assign M3nwx4 = (A4nwx4 & Lefwx4);
assign A4nwx4 = (~(H4nwx4 & W4zvx4));
assign W4zvx4 = (~(O4nwx4 & V4nwx4));
assign V4nwx4 = (C5nwx4 & J5nwx4);
assign J5nwx4 = (~(Wjyvx4 & Walwx4));
assign Wjyvx4 = (~(Q5nwx4 & X5nwx4));
assign X5nwx4 = (Iwdwx4 | E6nwx4);
assign Q5nwx4 = (~(L6nwx4 | S6nwx4));
assign L6nwx4 = (Z6nwx4 & G7nwx4);
assign Z6nwx4 = (~(N7nwx4 | Zph2z4[0]));
assign C5nwx4 = (U7nwx4 & Kkyvx4);
assign Kkyvx4 = (~(B8nwx4 & I8nwx4));
assign I8nwx4 = (~(P8nwx4 & W8nwx4));
assign P8nwx4 = (~(D9nwx4 & K9nwx4));
assign K9nwx4 = (Iwdwx4 & R9nwx4);
assign Iwdwx4 = (S1ewx4 | Y9nwx4);
assign D9nwx4 = (Fanwx4 & Z8ewx4);
assign Z8ewx4 = (~(Ay7wx4 & Manwx4));
assign U7nwx4 = (~(Amyvx4 & G9lwx4));
assign Amyvx4 = (~(Tanwx4 & Abnwx4));
assign Abnwx4 = (~(E6nwx4 & Hbnwx4));
assign Hbnwx4 = (~(Obnwx4 & Efgvx4));
assign Obnwx4 = (Vbnwx4 & Ccnwx4);
assign Ccnwx4 = (~(Jcnwx4 & Qcnwx4));
assign Qcnwx4 = (~(Dbgvx4 & Xcnwx4));
assign Xcnwx4 = (U9gvx4 | Mcgvx4);
assign Jcnwx4 = (~(Zph2z4[0] | Zph2z4[1]));
assign Vbnwx4 = (W5yvx4 | Bl3wx4);
assign O4nwx4 = (Ednwx4 & Ldnwx4);
assign Ldnwx4 = (~(Ykyvx4 & Palwx4));
assign Ykyvx4 = (~(Sdnwx4 & Zdnwx4));
assign Zdnwx4 = (~(Genwx4 & Ay7wx4));
assign Genwx4 = (Manwx4 & R9nwx4);
assign Sdnwx4 = (Nenwx4 & Uenwx4);
assign Nenwx4 = (~(Bfnwx4 & G7nwx4));
assign Bfnwx4 = (~(Ifnwx4 | N7nwx4));
assign Ednwx4 = (~(Omyvx4 & U9lwx4));
assign Omyvx4 = (~(Pfnwx4 & Wfnwx4));
assign Wfnwx4 = (Dgnwx4 & Kgnwx4);
assign Pfnwx4 = (~(Rgnwx4 | Ygnwx4));
assign Rgnwx4 = (Fhnwx4 & G7nwx4);
assign G7nwx4 = (Mhnwx4 & E6nwx4);
assign Mhnwx4 = (~(Dbgvx4 | Fjgvx4));
assign Fhnwx4 = (~(Ifnwx4 | Zph2z4[1]));
assign Y2nwx4 = (Thnwx4 & Ainwx4);
assign Ainwx4 = (~(Roh2z4[6] & Mifwx4));
assign Thnwx4 = (~(vis_pc_o[6] & Qaiwx4));
assign Skhvx4 = (~(Hinwx4 & Oinwx4));
assign Oinwx4 = (Vinwx4 & Cjnwx4);
assign Cjnwx4 = (~(Xdfwx4 & Dmh2z4[8]));
assign Vinwx4 = (Jjnwx4 & Lefwx4);
assign Jjnwx4 = (Sefwx4 | K22wx4);
assign K22wx4 = (Qjnwx4 & Xjnwx4);
assign Xjnwx4 = (Eknwx4 & Lknwx4);
assign Lknwx4 = (~(Sknwx4 & Hmyvx4));
assign Eknwx4 = (Zknwx4 & Glnwx4);
assign Zknwx4 = (~(Nlnwx4 & Pjyvx4));
assign Qjnwx4 = (Ulnwx4 & Bmnwx4);
assign Bmnwx4 = (~(Imnwx4 & Rkyvx4));
assign Ulnwx4 = (~(Pmnwx4 & Tlyvx4));
assign Hinwx4 = (Wmnwx4 & Dnnwx4);
assign Dnnwx4 = (~(Roh2z4[7] & Mifwx4));
assign Wmnwx4 = (~(vis_pc_o[7] & Qaiwx4));
assign Lkhvx4 = (~(Knnwx4 & Rnnwx4));
assign Rnnwx4 = (Ynnwx4 & Fonwx4);
assign Fonwx4 = (~(Xdfwx4 & Dmh2z4[10]));
assign Ynnwx4 = (Monwx4 & Lefwx4);
assign Monwx4 = (Sefwx4 | Wn1wx4);
assign Wn1wx4 = (Tonwx4 & Apnwx4);
assign Apnwx4 = (Hpnwx4 & Opnwx4);
assign Opnwx4 = (~(Nlnwx4 & Ajmwx4));
assign Hpnwx4 = (Vpnwx4 & Glnwx4);
assign Vpnwx4 = (~(Imnwx4 & Jkmwx4));
assign Tonwx4 = (Cqnwx4 & Jqnwx4);
assign Jqnwx4 = (~(Sknwx4 & Qkmwx4));
assign Cqnwx4 = (~(Pmnwx4 & Ojmwx4));
assign Knnwx4 = (Qqnwx4 & Xqnwx4);
assign Xqnwx4 = (~(Roh2z4[9] & Mifwx4));
assign Qqnwx4 = (~(vis_pc_o[9] & Qaiwx4));
assign Ekhvx4 = (~(Ernwx4 & Lrnwx4));
assign Lrnwx4 = (Srnwx4 & Zrnwx4);
assign Zrnwx4 = (~(Xdfwx4 & Dmh2z4[12]));
assign Srnwx4 = (Gsnwx4 & Lefwx4);
assign Gsnwx4 = (Sefwx4 | Uf1wx4);
assign Uf1wx4 = (Nsnwx4 & Usnwx4);
assign Usnwx4 = (Btnwx4 & Itnwx4);
assign Itnwx4 = (~(Sknwx4 & Xrmwx4));
assign Btnwx4 = (Ptnwx4 & Glnwx4);
assign Ptnwx4 = (~(Pmnwx4 & Gtmwx4));
assign Nsnwx4 = (Wtnwx4 & Dunwx4);
assign Dunwx4 = (~(Nlnwx4 & Ntmwx4));
assign Wtnwx4 = (~(Imnwx4 & Lsmwx4));
assign Ernwx4 = (Kunwx4 & Runwx4);
assign Runwx4 = (~(Roh2z4[11] & Mifwx4));
assign Kunwx4 = (~(vis_pc_o[11] & Qaiwx4));
assign Xjhvx4 = (~(Yunwx4 & Fvnwx4));
assign Fvnwx4 = (Mvnwx4 & Tvnwx4);
assign Tvnwx4 = (~(Xdfwx4 & Dmh2z4[14]));
assign Mvnwx4 = (Awnwx4 & Lefwx4);
assign Awnwx4 = (Sefwx4 | X61wx4);
assign X61wx4 = (Hwnwx4 & Ownwx4);
assign Ownwx4 = (Vwnwx4 & Cxnwx4);
assign Cxnwx4 = (~(Sknwx4 & D7iwx4));
assign Vwnwx4 = (Jxnwx4 & Glnwx4);
assign Jxnwx4 = (~(Nlnwx4 & Y7iwx4));
assign Hwnwx4 = (Qxnwx4 & Xxnwx4);
assign Xxnwx4 = (~(Imnwx4 & A9iwx4));
assign Qxnwx4 = (~(Pmnwx4 & O9iwx4));
assign Yunwx4 = (Eynwx4 & Lynwx4);
assign Lynwx4 = (~(Roh2z4[13] & Mifwx4));
assign Eynwx4 = (~(vis_pc_o[13] & Qaiwx4));
assign Qjhvx4 = (~(Synwx4 & Zynwx4));
assign Zynwx4 = (Gznwx4 & Nznwx4);
assign Nznwx4 = (~(Roh2z4[15] & Mifwx4));
assign Gznwx4 = (Uznwx4 & B0owx4);
assign B0owx4 = (Sefwx4 | I21wx4);
assign I21wx4 = (I0owx4 & P0owx4);
assign P0owx4 = (W0owx4 & D1owx4);
assign D1owx4 = (~(Yilwx4 & Pjyvx4));
assign Pjyvx4 = (~(K1owx4 & R1owx4));
assign R1owx4 = (Y1owx4 & F2owx4);
assign F2owx4 = (M2owx4 & T2owx4);
assign M2owx4 = (~(A3owx4 & Izgvx4));
assign A3owx4 = (A6tvx4 & H3owx4);
assign Y1owx4 = (O3owx4 & V3owx4);
assign V3owx4 = (~(W5rvx4 & C4owx4));
assign W5rvx4 = (J4owx4 & Q4owx4);
assign J4owx4 = (~(X4owx4 | E5owx4));
assign O3owx4 = (~(L5owx4 & U18wx4));
assign U18wx4 = (Yw7wx4 ? Xtdwx4 : E1ewx4);
assign K1owx4 = (S5owx4 & Z5owx4);
assign Z5owx4 = (~(Czh2z4[16] & G6owx4));
assign S5owx4 = (N6owx4 & U6owx4);
assign U6owx4 = (~(hrdata_i[16] & B7owx4));
assign N6owx4 = (~(Irh2z4[16] & I7owx4));
assign W0owx4 = (~(Phlwx4 & Hmyvx4));
assign Hmyvx4 = (~(P7owx4 & W7owx4));
assign W7owx4 = (D8owx4 & K8owx4);
assign K8owx4 = (~(L5owx4 & S08wx4));
assign S08wx4 = (Yw7wx4 ? C0ewx4 : Godwx4);
assign D8owx4 = (R8owx4 & Y8owx4);
assign Y8owx4 = (~(F9owx4 & L0i2z4[8]));
assign R8owx4 = (~(M9owx4 & T1i2z4[8]));
assign P7owx4 = (T9owx4 & Aaowx4);
assign Aaowx4 = (~(Czh2z4[8] & G6owx4));
assign T9owx4 = (Haowx4 & Oaowx4);
assign Oaowx4 = (~(hrdata_i[8] & B7owx4));
assign Haowx4 = (~(Irh2z4[8] & I7owx4));
assign I0owx4 = (Vaowx4 & Cbowx4);
assign Cbowx4 = (~(Fjlwx4 & Rkyvx4));
assign Rkyvx4 = (~(Jbowx4 & Qbowx4));
assign Qbowx4 = (~(hrdata_i[24] & B7owx4));
assign Jbowx4 = (Xbowx4 & Ecowx4);
assign Xbowx4 = (Lcowx4 | Q7ewx4);
assign Q7ewx4 = (Scowx4 & Zcowx4);
assign Zcowx4 = (Udowx4 ? Ndowx4 : Gdowx4);
assign Ndowx4 = (~(Yw7wx4 & Beowx4));
assign Gdowx4 = (Js7wx4 | M3ovx4);
assign Scowx4 = (Ieowx4 & Peowx4);
assign Peowx4 = (Weowx4 | Dfowx4);
assign Dfowx4 = (!Nvdwx4);
assign Ieowx4 = (~(Z08wx4 & M3ovx4));
assign Z08wx4 = (Yw7wx4 ? Beowx4 : Nvdwx4);
assign Vaowx4 = (~(W6iwx4 & Tlyvx4));
assign Tlyvx4 = (~(Kfowx4 & Rfowx4));
assign Rfowx4 = (Yfowx4 & Fgowx4);
assign Fgowx4 = (~(hrdata_i[0] & B7owx4));
assign Yfowx4 = (Mgowx4 & Tgowx4);
assign Tgowx4 = (~(H3owx4 & Ahowx4));
assign Ahowx4 = (~(Hhowx4 & Ohowx4));
assign Ohowx4 = (~(M5tvx4 & L0i2z4[0]));
assign Hhowx4 = (Vhowx4 & Ciowx4);
assign Ciowx4 = (~(F2hvx4 & A6tvx4));
assign Vhowx4 = (~(T1i2z4[0] & Ts5wx4));
assign Mgowx4 = (~(L5owx4 & B28wx4));
assign B28wx4 = (Yw7wx4 ? Qmdwx4 : Jiowx4);
assign Kfowx4 = (Qiowx4 & Xiowx4);
assign Xiowx4 = (~(Irh2z4[0] & I7owx4));
assign Qiowx4 = (~(Czh2z4[0] & G6owx4));
assign Uznwx4 = (~(Xdfwx4 & Dmh2z4[16]));
assign Synwx4 = (Tjlwx4 & Ejowx4);
assign Ejowx4 = (~(vis_pc_o[15] & Qaiwx4));
assign Jjhvx4 = (~(Ljowx4 & Sjowx4));
assign Sjowx4 = (Zjowx4 & Gkowx4);
assign Gkowx4 = (~(Roh2z4[16] & Mifwx4));
assign Zjowx4 = (Nkowx4 & Ukowx4);
assign Ukowx4 = (Sefwx4 | Mx0wx4);
assign Mx0wx4 = (Blowx4 & Ilowx4);
assign Ilowx4 = (Plowx4 & Wlowx4);
assign Wlowx4 = (~(W6iwx4 & Rhfwx4));
assign Plowx4 = (~(Phlwx4 & Khfwx4));
assign Blowx4 = (Dmowx4 & Kmowx4);
assign Kmowx4 = (~(Bgfwx4 & Yilwx4));
assign Dmowx4 = (~(Fjlwx4 & Pgfwx4));
assign Nkowx4 = (~(Xdfwx4 & Dmh2z4[17]));
assign Ljowx4 = (Tjlwx4 & Rmowx4);
assign Rmowx4 = (~(vis_pc_o[16] & Qaiwx4));
assign Cjhvx4 = (~(Ymowx4 & Fnowx4));
assign Fnowx4 = (Mnowx4 & Tnowx4);
assign Tnowx4 = (~(Roh2z4[17] & Mifwx4));
assign Mnowx4 = (Aoowx4 & Hoowx4);
assign Hoowx4 = (Sefwx4 | Et0wx4);
assign Et0wx4 = (Ooowx4 & Voowx4);
assign Voowx4 = (Cpowx4 & Jpowx4);
assign Jpowx4 = (~(Fjlwx4 & Jkmwx4));
assign Cpowx4 = (~(Ajmwx4 & Yilwx4));
assign Ooowx4 = (Qpowx4 & Xpowx4);
assign Xpowx4 = (~(Phlwx4 & Qkmwx4));
assign Qpowx4 = (~(W6iwx4 & Ojmwx4));
assign Aoowx4 = (~(Xdfwx4 & Dmh2z4[18]));
assign Ymowx4 = (Tjlwx4 & Eqowx4);
assign Eqowx4 = (~(vis_pc_o[17] & Qaiwx4));
assign Vihvx4 = (~(Lqowx4 & Sqowx4));
assign Sqowx4 = (Zqowx4 & Growx4);
assign Growx4 = (~(Roh2z4[21] & Mifwx4));
assign Zqowx4 = (Nrowx4 & Urowx4);
assign Urowx4 = (Sefwx4 | Ba0wx4);
assign Ba0wx4 = (Bsowx4 & Isowx4);
assign Isowx4 = (Psowx4 & Wsowx4);
assign Wsowx4 = (~(Y7iwx4 & Yilwx4));
assign Y7iwx4 = (~(Dtowx4 & Ktowx4));
assign Ktowx4 = (Rtowx4 & Ytowx4);
assign Ytowx4 = (~(Fuowx4 & Muowx4));
assign Rtowx4 = (Tuowx4 & Avowx4);
assign Avowx4 = (~(H3owx4 & Hvowx4));
assign Hvowx4 = (~(Ovowx4 & Vvowx4));
assign Vvowx4 = (Cwowx4 & Jwowx4);
assign Jwowx4 = (Qwowx4 | Xwowx4);
assign Cwowx4 = (Exowx4 & Lxowx4);
assign Lxowx4 = (K3uvx4 | Sxowx4);
assign Exowx4 = (E0uvx4 | Zxowx4);
assign Ovowx4 = (Gyowx4 & Nyowx4);
assign Nyowx4 = (~(S0uvx4 & Zuh2z4[12]));
assign Gyowx4 = (N1uvx4 | Uyowx4);
assign Tuowx4 = (~(Bzowx4 & Zudwx4));
assign Dtowx4 = (Izowx4 & Pzowx4);
assign Pzowx4 = (~(Czh2z4[22] & G6owx4));
assign Izowx4 = (Wzowx4 & D0pwx4);
assign D0pwx4 = (~(hrdata_i[22] & B7owx4));
assign Wzowx4 = (~(Irh2z4[22] & I7owx4));
assign Psowx4 = (~(Phlwx4 & D7iwx4));
assign D7iwx4 = (~(K0pwx4 & R0pwx4));
assign R0pwx4 = (Y0pwx4 & F1pwx4);
assign F1pwx4 = (~(H3owx4 & M1pwx4));
assign M1pwx4 = (~(T1pwx4 & A2pwx4));
assign A2pwx4 = (H2pwx4 & O2pwx4);
assign O2pwx4 = (V2pwx4 & C3pwx4);
assign C3pwx4 = (E0uvx4 | J3pwx4);
assign V2pwx4 = (Q3pwx4 & X3pwx4);
assign Q3pwx4 = (~(X2rvx4 & Gc4wx4));
assign X2rvx4 = (~(E4pwx4 | L4pwx4));
assign E4pwx4 = (G5pwx4 ? Z4pwx4 : S4pwx4);
assign Z4pwx4 = (~(X4owx4 | N5pwx4));
assign N5pwx4 = (I6pwx4 ? B6pwx4 : U5pwx4);
assign H2pwx4 = (P6pwx4 & W6pwx4);
assign W6pwx4 = (Qwowx4 | D7pwx4);
assign P6pwx4 = (K7pwx4 | R7pwx4);
assign T1pwx4 = (Y7pwx4 & F8pwx4);
assign F8pwx4 = (M8pwx4 & T8pwx4);
assign T8pwx4 = (~(M5tvx4 & L0i2z4[14]));
assign M8pwx4 = (A9pwx4 & H9pwx4);
assign H9pwx4 = (N1uvx4 | O9pwx4);
assign A9pwx4 = (~(T1i2z4[14] & Ts5wx4));
assign Y7pwx4 = (V9pwx4 & Capwx4);
assign Capwx4 = (~(Irh2z4[14] & Japwx4));
assign V9pwx4 = (~(Czh2z4[14] & H6tvx4));
assign Y0pwx4 = (~(Bzowx4 & Eudwx4));
assign K0pwx4 = (Qapwx4 & Xapwx4);
assign Xapwx4 = (~(Fuowx4 & Ebpwx4));
assign Qapwx4 = (~(hrdata_i[14] & B7owx4));
assign Bsowx4 = (Lbpwx4 & Sbpwx4);
assign Sbpwx4 = (~(Fjlwx4 & A9iwx4));
assign A9iwx4 = (~(Zbpwx4 & Gcpwx4));
assign Gcpwx4 = (~(hrdata_i[30] & B7owx4));
assign Zbpwx4 = (Ncpwx4 & Ucpwx4);
assign Ucpwx4 = (~(L5owx4 & J7ewx4));
assign J7ewx4 = (Idpwx4 ? U2ewx4 : Bdpwx4);
assign Idpwx4 = (Pdpwx4 & Wdpwx4);
assign Pdpwx4 = (Depwx4 ? Weowx4 : Udowx4);
assign Bdpwx4 = (Oldwx4 ? Kepwx4 : Xmdwx4);
assign Ncpwx4 = (~(H3owx4 & Repwx4));
assign Repwx4 = (~(Yepwx4 & Ffpwx4));
assign Ffpwx4 = (Mfpwx4 & Tfpwx4);
assign Tfpwx4 = (Agpwx4 & X3pwx4);
assign Agpwx4 = (~(P2uvx4 & Uth2z4[0]));
assign Mfpwx4 = (Hgpwx4 & Ogpwx4);
assign Ogpwx4 = (K3uvx4 | Vgpwx4);
assign Hgpwx4 = (E0uvx4 | Chpwx4);
assign Yepwx4 = (Jhpwx4 & Qhpwx4);
assign Qhpwx4 = (Xhpwx4 & Eipwx4);
assign Eipwx4 = (Qwowx4 | Lipwx4);
assign Xhpwx4 = (K7pwx4 | Sipwx4);
assign Jhpwx4 = (Zipwx4 & Gjpwx4);
assign Gjpwx4 = (N1uvx4 | Njpwx4);
assign Lbpwx4 = (~(W6iwx4 & O9iwx4));
assign O9iwx4 = (~(Ujpwx4 & Bkpwx4));
assign Bkpwx4 = (Ikpwx4 & Pkpwx4);
assign Pkpwx4 = (~(H3owx4 & Wkpwx4));
assign Wkpwx4 = (~(Dlpwx4 & Klpwx4));
assign Klpwx4 = (Rlpwx4 & Ylpwx4);
assign Ylpwx4 = (Fmpwx4 & Mmpwx4);
assign Mmpwx4 = (E0uvx4 | Tmpwx4);
assign Fmpwx4 = (~(Jztvx4 & Zuh2z4[24]));
assign Jztvx4 = (!Qwowx4);
assign Rlpwx4 = (Anpwx4 & Hnpwx4);
assign Hnpwx4 = (~(S0uvx4 & Zuh2z4[8]));
assign S0uvx4 = (!K7pwx4);
assign Anpwx4 = (N1uvx4 | Onpwx4);
assign Dlpwx4 = (Vnpwx4 & Copwx4);
assign Copwx4 = (Jopwx4 & Qopwx4);
assign Qopwx4 = (~(T1i2z4[6] & Ts5wx4));
assign Jopwx4 = (~(M5tvx4 & L0i2z4[6]));
assign Vnpwx4 = (Xopwx4 & Eppwx4);
assign Eppwx4 = (~(Irh2z4[6] & Japwx4));
assign Xopwx4 = (~(Czh2z4[6] & H6tvx4));
assign Ikpwx4 = (~(Bzowx4 & Sndwx4));
assign Ujpwx4 = (Lppwx4 & Sppwx4);
assign Sppwx4 = (~(Fuowx4 & Zppwx4));
assign Lppwx4 = (~(hrdata_i[6] & B7owx4));
assign Nrowx4 = (~(Xdfwx4 & Dmh2z4[22]));
assign Lqowx4 = (Tjlwx4 & Gqpwx4);
assign Gqpwx4 = (~(vis_pc_o[21] & Qaiwx4));
assign Oihvx4 = (~(Nqpwx4 & Uqpwx4));
assign Uqpwx4 = (Brpwx4 & Irpwx4);
assign Irpwx4 = (~(Xdfwx4 & Dmh2z4[25]));
assign Brpwx4 = (Prpwx4 & Lefwx4);
assign Prpwx4 = (Sefwx4 | Ppzvx4);
assign Ppzvx4 = (Wrpwx4 & Dspwx4);
assign Dspwx4 = (Kspwx4 & Rspwx4);
assign Rspwx4 = (~(Rhfwx4 & V9iwx4));
assign Kspwx4 = (Yspwx4 & R7iwx4);
assign Yspwx4 = (~(Pgfwx4 & H9iwx4));
assign Wrpwx4 = (Ftpwx4 & Mtpwx4);
assign Mtpwx4 = (~(W6iwx4 & Khfwx4));
assign Ftpwx4 = (~(Bgfwx4 & F8iwx4));
assign Nqpwx4 = (Ttpwx4 & Aupwx4);
assign Aupwx4 = (~(Roh2z4[24] & Mifwx4));
assign Ttpwx4 = (~(vis_pc_o[24] & Qaiwx4));
assign Hihvx4 = (~(Hupwx4 & Oupwx4));
assign Oupwx4 = (Vupwx4 & Cvpwx4);
assign Cvpwx4 = (~(Xdfwx4 & Dmh2z4[26]));
assign Vupwx4 = (Jvpwx4 & Lefwx4);
assign Jvpwx4 = (Sefwx4 | Yjzvx4);
assign Yjzvx4 = (Qvpwx4 & Xvpwx4);
assign Xvpwx4 = (Ewpwx4 & Lwpwx4);
assign Lwpwx4 = (~(Ajmwx4 & F8iwx4));
assign Ajmwx4 = (~(Swpwx4 & Zwpwx4));
assign Zwpwx4 = (Gxpwx4 & Nxpwx4);
assign Nxpwx4 = (T2owx4 & Ecowx4);
assign Gxpwx4 = (Uxpwx4 & Bypwx4);
assign Bypwx4 = (~(Fuowx4 & Eudwx4));
assign Eudwx4 = (~(Iypwx4 & Pypwx4));
assign Pypwx4 = (Wypwx4 & Dzpwx4);
assign Dzpwx4 = (~(Kzpwx4 & Rzpwx4));
assign Wypwx4 = (~(Yzpwx4 & F0qwx4));
assign Iypwx4 = (M0qwx4 & T0qwx4);
assign T0qwx4 = (A1qwx4 | H1qwx4);
assign M0qwx4 = (~(O1qwx4 & V1qwx4));
assign Uxpwx4 = (~(Bzowx4 & Muowx4));
assign Muowx4 = (!Asdwx4);
assign Asdwx4 = (C2qwx4 & J2qwx4);
assign J2qwx4 = (Q2qwx4 & X2qwx4);
assign X2qwx4 = (~(Kzpwx4 & E3qwx4));
assign Q2qwx4 = (~(O1qwx4 & L3qwx4));
assign C2qwx4 = (S3qwx4 & Z3qwx4);
assign Z3qwx4 = (A1qwx4 | G4qwx4);
assign S3qwx4 = (~(Yzpwx4 & N4qwx4));
assign Swpwx4 = (U4qwx4 & B5qwx4);
assign B5qwx4 = (~(Czh2z4[18] & G6owx4));
assign U4qwx4 = (I5qwx4 & P5qwx4);
assign P5qwx4 = (~(hrdata_i[18] & B7owx4));
assign I5qwx4 = (~(Irh2z4[18] & I7owx4));
assign Ewpwx4 = (W5qwx4 & R7iwx4);
assign W5qwx4 = (~(Jkmwx4 & H9iwx4));
assign Jkmwx4 = (~(D6qwx4 & K6qwx4));
assign K6qwx4 = (R6qwx4 & Y6qwx4);
assign Y6qwx4 = (F7qwx4 | M7qwx4);
assign R6qwx4 = (~(C4owx4 & R3hvx4));
assign D6qwx4 = (T7qwx4 & A8qwx4);
assign A8qwx4 = (A6ewx4 | Lcowx4);
assign A6ewx4 = (~(H8qwx4 & F7qwx4));
assign F7qwx4 = (O8qwx4 | V8qwx4);
assign O8qwx4 = (Depwx4 ? Udowx4 : C9qwx4);
assign H8qwx4 = (Yw7wx4 ? Kepwx4 : Zudwx4);
assign Kepwx4 = (~(J9qwx4 & Q9qwx4));
assign Q9qwx4 = (X9qwx4 & Eaqwx4);
assign Eaqwx4 = (~(O1qwx4 & Laqwx4));
assign X9qwx4 = (A1qwx4 | Saqwx4);
assign J9qwx4 = (Zaqwx4 & Gbqwx4);
assign Gbqwx4 = (~(Yzpwx4 & Nbqwx4));
assign Zaqwx4 = (~(Kzpwx4 & Ubqwx4));
assign Zudwx4 = (~(Bcqwx4 & Icqwx4));
assign Icqwx4 = (Pcqwx4 & Wcqwx4);
assign Wcqwx4 = (~(Kzpwx4 & Ddqwx4));
assign Pcqwx4 = (~(Yzpwx4 & Kdqwx4));
assign Bcqwx4 = (Rdqwx4 & Ydqwx4);
assign Ydqwx4 = (A1qwx4 | Feqwx4);
assign Rdqwx4 = (~(O1qwx4 & Meqwx4));
assign T7qwx4 = (~(hrdata_i[26] & B7owx4));
assign Qvpwx4 = (Teqwx4 & Afqwx4);
assign Afqwx4 = (~(W6iwx4 & Qkmwx4));
assign Qkmwx4 = (~(Hfqwx4 & Ofqwx4));
assign Ofqwx4 = (Vfqwx4 & Cgqwx4);
assign Cgqwx4 = (Jgqwx4 & Qgqwx4);
assign Qgqwx4 = (~(F9owx4 & L0i2z4[10]));
assign Jgqwx4 = (~(M9owx4 & T1i2z4[10]));
assign Vfqwx4 = (Xgqwx4 & Ehqwx4);
assign Ehqwx4 = (~(Fuowx4 & Sndwx4));
assign Sndwx4 = (~(Lhqwx4 & Shqwx4));
assign Shqwx4 = (Zhqwx4 & Giqwx4);
assign Giqwx4 = (~(Kzpwx4 & Niqwx4));
assign Zhqwx4 = (~(Yzpwx4 & Uiqwx4));
assign Lhqwx4 = (Bjqwx4 & Ijqwx4);
assign Ijqwx4 = (A1qwx4 | Pjqwx4);
assign Bjqwx4 = (~(O1qwx4 & Wjqwx4));
assign Xgqwx4 = (~(Bzowx4 & Ebpwx4));
assign Ebpwx4 = (!Mydwx4);
assign Mydwx4 = (Dkqwx4 & Kkqwx4);
assign Kkqwx4 = (Rkqwx4 & Ykqwx4);
assign Ykqwx4 = (~(Kzpwx4 & Flqwx4));
assign Rkqwx4 = (~(O1qwx4 & Mlqwx4));
assign Dkqwx4 = (Tlqwx4 & Amqwx4);
assign Amqwx4 = (A1qwx4 | Hmqwx4);
assign Tlqwx4 = (~(Yzpwx4 & Omqwx4));
assign Hfqwx4 = (Vmqwx4 & Cnqwx4);
assign Cnqwx4 = (~(Czh2z4[10] & G6owx4));
assign Vmqwx4 = (Jnqwx4 & Qnqwx4);
assign Qnqwx4 = (~(hrdata_i[10] & B7owx4));
assign Jnqwx4 = (~(Irh2z4[10] & I7owx4));
assign Teqwx4 = (~(Ojmwx4 & V9iwx4));
assign Ojmwx4 = (~(Xnqwx4 & Eoqwx4));
assign Eoqwx4 = (Loqwx4 & Soqwx4);
assign Soqwx4 = (~(Fuowx4 & Xmdwx4));
assign Xmdwx4 = (~(Zoqwx4 & Gpqwx4));
assign Gpqwx4 = (Npqwx4 & Upqwx4);
assign Upqwx4 = (~(Kzpwx4 & Bqqwx4));
assign Npqwx4 = (~(Yzpwx4 & Iqqwx4));
assign Zoqwx4 = (Pqqwx4 & Wqqwx4);
assign Wqqwx4 = (A1qwx4 | Ylbwx4);
assign Pqqwx4 = (~(O1qwx4 & Drqwx4));
assign Loqwx4 = (Krqwx4 & Rrqwx4);
assign Rrqwx4 = (~(H3owx4 & Yrqwx4));
assign Yrqwx4 = (~(Fsqwx4 & Msqwx4));
assign Msqwx4 = (Tsqwx4 & A5uvx4);
assign Tsqwx4 = (~(T1i2z4[2] & Ts5wx4));
assign Fsqwx4 = (Atqwx4 & Htqwx4);
assign Htqwx4 = (~(Nngvx4 & B2uvx4));
assign Atqwx4 = (~(M5tvx4 & L0i2z4[2]));
assign Krqwx4 = (~(Bzowx4 & Zppwx4));
assign Zppwx4 = (!Tkdwx4);
assign Tkdwx4 = (Otqwx4 & Vtqwx4);
assign Vtqwx4 = (Cuqwx4 & Juqwx4);
assign Juqwx4 = (~(Kzpwx4 & Quqwx4));
assign Cuqwx4 = (~(O1qwx4 & Xuqwx4));
assign Otqwx4 = (Evqwx4 & Lvqwx4);
assign Lvqwx4 = (A1qwx4 | Svqwx4);
assign Evqwx4 = (~(Yzpwx4 & Zvqwx4));
assign Xnqwx4 = (Gwqwx4 & Nwqwx4);
assign Nwqwx4 = (~(Czh2z4[2] & G6owx4));
assign Gwqwx4 = (Uwqwx4 & Bxqwx4);
assign Bxqwx4 = (~(hrdata_i[2] & B7owx4));
assign Uwqwx4 = (~(Irh2z4[2] & I7owx4));
assign Hupwx4 = (Ixqwx4 & Pxqwx4);
assign Pxqwx4 = (~(Roh2z4[25] & Mifwx4));
assign Ixqwx4 = (~(vis_pc_o[25] & Qaiwx4));
assign Aihvx4 = (~(Wxqwx4 & Dyqwx4));
assign Dyqwx4 = (Kyqwx4 & Ryqwx4);
assign Ryqwx4 = (~(Xdfwx4 & Dmh2z4[27]));
assign Kyqwx4 = (Yyqwx4 & Lefwx4);
assign Yyqwx4 = (Sefwx4 | Qfzvx4);
assign Qfzvx4 = (Fzqwx4 & Mzqwx4);
assign Mzqwx4 = (Tzqwx4 & A0rwx4);
assign A0rwx4 = (~(Ihlwx4 & V9iwx4));
assign Tzqwx4 = (H0rwx4 & R7iwx4);
assign H0rwx4 = (~(Mjlwx4 & H9iwx4));
assign Fzqwx4 = (O0rwx4 & V0rwx4);
assign V0rwx4 = (~(W6iwx4 & Whlwx4));
assign O0rwx4 = (~(Rilwx4 & F8iwx4));
assign Wxqwx4 = (C1rwx4 & J1rwx4);
assign J1rwx4 = (~(Roh2z4[26] & Mifwx4));
assign C1rwx4 = (~(vis_pc_o[26] & Qaiwx4));
assign Thhvx4 = (~(Q1rwx4 & X1rwx4));
assign X1rwx4 = (E2rwx4 & L2rwx4);
assign L2rwx4 = (~(Xdfwx4 & Dmh2z4[28]));
assign E2rwx4 = (S2rwx4 & Lefwx4);
assign S2rwx4 = (Sefwx4 | Wzpvx4);
assign Wzpvx4 = (Z2rwx4 & G3rwx4);
assign G3rwx4 = (N3rwx4 & U3rwx4);
assign U3rwx4 = (~(Lsmwx4 & H9iwx4));
assign N3rwx4 = (B4rwx4 & R7iwx4);
assign B4rwx4 = (~(W6iwx4 & Xrmwx4));
assign Z2rwx4 = (I4rwx4 & P4rwx4);
assign P4rwx4 = (~(Gtmwx4 & V9iwx4));
assign I4rwx4 = (~(Ntmwx4 & F8iwx4));
assign Q1rwx4 = (W4rwx4 & D5rwx4);
assign D5rwx4 = (~(Roh2z4[27] & Mifwx4));
assign W4rwx4 = (~(vis_pc_o[27] & Qaiwx4));
assign Mhhvx4 = (~(K5rwx4 & R5rwx4));
assign R5rwx4 = (Y5rwx4 & F6rwx4);
assign F6rwx4 = (~(Xdfwx4 & Dmh2z4[29]));
assign Y5rwx4 = (M6rwx4 & Lefwx4);
assign M6rwx4 = (Sefwx4 | Bspvx4);
assign Bspvx4 = (T6rwx4 & A7rwx4);
assign A7rwx4 = (H7rwx4 & O7rwx4);
assign O7rwx4 = (~(Cymwx4 & V9iwx4));
assign V9iwx4 = (~(Uenwx4 & V7rwx4));
assign V7rwx4 = (C8rwx4 | Z1ewx4);
assign H7rwx4 = (J8rwx4 & R7iwx4);
assign R7iwx4 = (~(Q8rwx4 & X8rwx4));
assign X8rwx4 = (~(Cs7wx4 & R9nwx4));
assign Cs7wx4 = (~(E9rwx4 & Ipdwx4));
assign Ipdwx4 = (~(Dp7wx4 & L9rwx4));
assign L9rwx4 = (Mq7wx4 | Yp7wx4);
assign E9rwx4 = (Qs7wx4 & S8ewx4);
assign J8rwx4 = (~(Hxmwx4 & H9iwx4));
assign H9iwx4 = (~(S9rwx4 & Z9rwx4));
assign Z9rwx4 = (S8ewx4 | E6nwx4);
assign T6rwx4 = (Garwx4 & Narwx4);
assign Narwx4 = (~(Jymwx4 & F8iwx4));
assign Garwx4 = (~(W6iwx4 & Twmwx4));
assign K5rwx4 = (Uarwx4 & Bbrwx4);
assign Bbrwx4 = (~(Roh2z4[28] & Mifwx4));
assign Uarwx4 = (~(vis_pc_o[28] & Qaiwx4));
assign Fhhvx4 = (hready_i ? Ibrwx4 : A3gvx4);
assign Ibrwx4 = (~(Pbrwx4 & Wbrwx4));
assign Wbrwx4 = (Dcrwx4 | A3gvx4);
assign Pbrwx4 = (Kcrwx4 & Rcrwx4);
assign Rcrwx4 = (Y8pvx4 | Hlsvx4);
assign Kcrwx4 = (~(I4gvx4 & Ipsvx4));
assign Yghvx4 = (~(Ycrwx4 & Fdrwx4));
assign Fdrwx4 = (~(Mdrwx4 & A3gvx4));
assign Mdrwx4 = (Tdrwx4 & hready_i);
assign Tdrwx4 = (~(Dcrwx4 & S5pvx4));
assign Ycrwx4 = (~(I4gvx4 & Aerwx4));
assign Aerwx4 = (~(G6pvx4 & S5pvx4));
assign Rghvx4 = (Yafwx4 ? Herwx4 : Tjh2z4[2]);
assign Yafwx4 = (Oerwx4 & hready_i);
assign Oerwx4 = (~(Verwx4 & Cfrwx4));
assign Cfrwx4 = (Jfrwx4 & Qfrwx4);
assign Qfrwx4 = (~(Xfrwx4 & M1xvx4));
assign Xfrwx4 = (~(Egrwx4 & Lgrwx4));
assign Lgrwx4 = (Sgrwx4 & Zgrwx4);
assign Zgrwx4 = (~(Ghrwx4 & Cn8vx4));
assign Ghrwx4 = (Nhrwx4 & Lcpvx4);
assign Nhrwx4 = (~(Oigwx4 & Y5svx4));
assign Oigwx4 = (Qfsvx4 & Dfpvx4);
assign Sgrwx4 = (~(Ovwvx4 | Mk6wx4));
assign Ovwvx4 = (Wi6wx4 & Q4wvx4);
assign Q4wvx4 = (~(Bisvx4 | Izwvx4));
assign Wi6wx4 = (~(Xmsvx4 | Ud9vx4));
assign Egrwx4 = (Uhrwx4 & Birwx4);
assign Birwx4 = (~(Xhxvx4 & Iirwx4));
assign Iirwx4 = (Abgwx4 | Xmsvx4);
assign Uhrwx4 = (Dziwx4 | Y99vx4);
assign Jfrwx4 = (~(Pirwx4 | Cp3wx4));
assign Cp3wx4 = (~(Dziwx4 | Lcpvx4));
assign Dziwx4 = (!Nkpvx4);
assign Pirwx4 = (Wirwx4 & Lxwvx4);
assign Wirwx4 = (~(Mc9vx4 | Y99vx4));
assign Verwx4 = (Djrwx4 & J3xvx4);
assign J3xvx4 = (Kjrwx4 & Rjrwx4);
assign Rjrwx4 = (~(Wshwx4 & Yjrwx4));
assign Yjrwx4 = (~(Ct6wx4 & Fkrwx4));
assign Fkrwx4 = (~(A4gwx4 & J16wx4));
assign A4gwx4 = (~(Lqwvx4 | Y99vx4));
assign Wshwx4 = (!Qoiwx4);
assign Kjrwx4 = (~(Mkrwx4 | Mljwx4));
assign Djrwx4 = (Tkrwx4 & Alrwx4);
assign Alrwx4 = (Sznvx4 | F57wx4);
assign Tkrwx4 = (Gjxvx4 | Whgvx4);
assign Gjxvx4 = (!M66wx4);
assign Herwx4 = (~(Hlrwx4 & Olrwx4));
assign Olrwx4 = (Vlrwx4 & Cmrwx4);
assign Cmrwx4 = (Fdsvx4 | J3iwx4);
assign J3iwx4 = (Lcpvx4 ? Qmrwx4 : Jmrwx4);
assign Qmrwx4 = (~(Xmrwx4 & Kg9vx4));
assign Xmrwx4 = (~(U4yvx4 | Sh9vx4));
assign Vlrwx4 = (~(Q3iwx4 & D69vx4));
assign Q3iwx4 = (Rngwx4 & Enrwx4);
assign Enrwx4 = (~(Lnrwx4 & Dthwx4));
assign Dthwx4 = (!Qsewx4);
assign Lnrwx4 = (Dfpvx4 ? Znrwx4 : Snrwx4);
assign Znrwx4 = (Cf9vx4 ? Aj9vx4 : Sh9vx4);
assign Snrwx4 = (Epxvx4 | Uasvx4);
assign Hlrwx4 = (Fbfwx4 & Gorwx4);
assign Gorwx4 = (~(I29vx4 & E4iwx4));
assign E4iwx4 = (~(Ocfwx4 & Norwx4));
assign Norwx4 = (Acfwx4 | P39vx4);
assign Fbfwx4 = (Uorwx4 & Bprwx4);
assign Bprwx4 = (Iprwx4 & Pprwx4);
assign Pprwx4 = (~(Fjgvx4 & Wprwx4));
assign Wprwx4 = (M3ovx4 | P39vx4);
assign Iprwx4 = (Dqrwx4 & Bswvx4);
assign Bswvx4 = (!Fv2wx4);
assign Dqrwx4 = (~(Jjgwx4 & Kqrwx4));
assign Kqrwx4 = (Uasvx4 | Dfpvx4);
assign Uorwx4 = (Celwx4 & Rqrwx4);
assign Rqrwx4 = (~(Kg9vx4 & K8hwx4));
assign Celwx4 = (Yqrwx4 & Frrwx4);
assign Frrwx4 = (Ocfwx4 | Mrrwx4);
assign Mrrwx4 = (Qfsvx4 & Trrwx4);
assign Trrwx4 = (Abgwx4 | J8svx4);
assign Ocfwx4 = (~(Asrwx4 & Hsrwx4));
assign Hsrwx4 = (~(Kg9vx4 | Aj9vx4));
assign Asrwx4 = (~(Jmrwx4 | Cf9vx4));
assign Yqrwx4 = (~(Osrwx4 | Keiwx4));
assign Keiwx4 = (~(Jmrwx4 | Epxvx4));
assign Jmrwx4 = (Xmsvx4 | U4yvx4);
assign Osrwx4 = (Vsrwx4 & Nakwx4);
assign Nakwx4 = (~(Uz8vx4 | B19vx4));
assign Vsrwx4 = (~(Gwrvx4 | Acfwx4));
assign Kghvx4 = (~(Ctrwx4 & Jtrwx4));
assign Jtrwx4 = (~(Qtrwx4 & Cllwx4));
assign Ctrwx4 = (Qllwx4 ? Xtrwx4 : Cwawx4);
assign Xtrwx4 = (Eurwx4 & Lurwx4);
assign Lurwx4 = (Surwx4 & Zurwx4);
assign Zurwx4 = (~(Orlwx4 & Fuevx4));
assign Orlwx4 = (~(Wyxvx4 | Gvrwx4));
assign Gvrwx4 = (Nvrwx4 & Vp2wx4);
assign Nvrwx4 = (~(Uvrwx4 | P5yvx4));
assign Wyxvx4 = (!Xlevx4);
assign Surwx4 = (~(D69vx4 & Vrlwx4));
assign Eurwx4 = (Bwrwx4 & Iwrwx4);
assign Iwrwx4 = (~(Dsqvx4 & Mc9vx4));
assign Dsqvx4 = (Mljwx4 & C2yvx4);
assign Bwrwx4 = (~(W49vx4 & Qslwx4));
assign Dghvx4 = (Pwrwx4 | Wwrwx4);
assign Wwrwx4 = (Dxrwx4 & Cllwx4);
assign Pwrwx4 = (Qllwx4 ? Kxrwx4 : Gr9vx4);
assign Kxrwx4 = (~(Rxrwx4 & Yxrwx4));
assign Yxrwx4 = (~(K79vx4 & Vrlwx4));
assign Vrlwx4 = (Fyrwx4 | Ohwvx4);
assign Rxrwx4 = (~(D69vx4 & Qslwx4));
assign Wfhvx4 = (Myrwx4 | Tyrwx4);
assign Tyrwx4 = (Azrwx4 & Cllwx4);
assign Cllwx4 = (~(Hzrwx4 & Dplwx4));
assign Dplwx4 = (Ozrwx4 & Vzrwx4);
assign Vzrwx4 = (Sznvx4 | Xviwx4);
assign Ozrwx4 = (Lbiwx4 | Nggvx4);
assign Hzrwx4 = (C0swx4 & Arewx4);
assign Arewx4 = (!Agbwx4);
assign Agbwx4 = (Fjgvx4 & U9gvx4);
assign C0swx4 = (~(C9yvx4 & Rngwx4));
assign Myrwx4 = (Qllwx4 ? J0swx4 : Ks9vx4);
assign Qllwx4 = (Q0swx4 & hready_i);
assign Q0swx4 = (~(X0swx4 & E1swx4));
assign E1swx4 = (L1swx4 & S1swx4);
assign S1swx4 = (Z1swx4 & G2swx4);
assign G2swx4 = (~(N2swx4 & Q5gvx4));
assign N2swx4 = (Pkxvx4 & Huqvx4);
assign Z1swx4 = (~(Wdxvx4 & Jwwvx4));
assign L1swx4 = (U2swx4 & B3swx4);
assign B3swx4 = (~(I3swx4 & B1vvx4));
assign U2swx4 = (Qoiwx4 | Kg9vx4);
assign X0swx4 = (P3swx4 & Q3xvx4);
assign Q3xvx4 = (W3swx4 & D4swx4);
assign D4swx4 = (~(D13wx4 & W9fwx4));
assign W3swx4 = (K4swx4 & R4swx4);
assign R4swx4 = (~(Y4swx4 & A0zvx4));
assign Y4swx4 = (~(U9gvx4 | Mcgvx4));
assign K4swx4 = (Jhxvx4 | Wqjwx4);
assign Wqjwx4 = (!Pa7wx4);
assign P3swx4 = (Bkxvx4 & F5swx4);
assign F5swx4 = (~(M5swx4 & Ju5wx4));
assign Bkxvx4 = (T5swx4 & A6swx4);
assign A6swx4 = (H6swx4 & O6swx4);
assign O6swx4 = (Ae6wx4 & Lbiwx4);
assign Ae6wx4 = (~(V6swx4 & Izwvx4));
assign H6swx4 = (C7swx4 & J7swx4);
assign J7swx4 = (~(Lxwvx4 & Q7swx4));
assign Q7swx4 = (Sh9vx4 | Tr6wx4);
assign Tr6wx4 = (~(Y99vx4 | Fb9vx4));
assign Lxwvx4 = (!H5fwx4);
assign H5fwx4 = (~(Wvewx4 & Qfsvx4));
assign C7swx4 = (Ct6wx4 | Qoiwx4);
assign Qoiwx4 = (~(Wvewx4 & Xmsvx4));
assign Ct6wx4 = (!Ksiwx4);
assign Ksiwx4 = (~(Fdsvx4 | Fb9vx4));
assign T5swx4 = (X7swx4 & E8swx4);
assign E8swx4 = (L8swx4 & S8swx4);
assign S8swx4 = (~(Z8swx4 & M1xvx4));
assign Z8swx4 = (~(G9swx4 & N9swx4));
assign N9swx4 = (~(U9swx4 | Nzgwx4));
assign U9swx4 = (Nkpvx4 & Baswx4);
assign Baswx4 = (~(Iaswx4 & Paswx4));
assign Paswx4 = (~(Dj6wx4 & H4gwx4));
assign H4gwx4 = (Y99vx4 & Zn6wx4);
assign Iaswx4 = (Abgwx4 | Fk6wx4);
assign Fk6wx4 = (!Uijwx4);
assign Uijwx4 = (~(J8svx4 | Y5svx4));
assign Nkpvx4 = (~(Iufwx4 | Ud9vx4));
assign G9swx4 = (Waswx4 & Dbswx4);
assign Dbswx4 = (X5gwx4 | Sh9vx4);
assign Waswx4 = (Yj6wx4 | Aj9vx4);
assign L8swx4 = (Fzyvx4 | P39vx4);
assign X7swx4 = (X3xvx4 & Bw6wx4);
assign Bw6wx4 = (Svyvx4 & Kbswx4);
assign Kbswx4 = (~(T1xvx4 & W5yvx4));
assign Svyvx4 = (!Mkrwx4);
assign Mkrwx4 = (Fv2wx4 & Z2zvx4);
assign Z2zvx4 = (!Msyvx4);
assign Fv2wx4 = (~(O4ovx4 | Fjgvx4));
assign X3xvx4 = (Rbswx4 & Ybswx4);
assign Ybswx4 = (Fcswx4 & Eqhwx4);
assign Eqhwx4 = (Ulgwx4 | Lcpvx4);
assign Ulgwx4 = (!Mk6wx4);
assign Mk6wx4 = (~(Iufwx4 | Sh9vx4));
assign Fcswx4 = (~(Mcswx4 & Wvewx4));
assign Mcswx4 = (~(G27wx4 | Kg9vx4));
assign Rbswx4 = (Tcswx4 & Adswx4);
assign Adswx4 = (~(Hdswx4 & Eznvx4));
assign Hdswx4 = (~(H33wx4 | Cn8vx4));
assign Tcswx4 = (Fzyvx4 | U9gvx4);
assign Fzyvx4 = (~(Srgwx4 & Zrvvx4));
assign J0swx4 = (~(Odswx4 & Vdswx4));
assign Vdswx4 = (~(R89vx4 & Fyrwx4));
assign Fyrwx4 = (~(Ceswx4 & Jeswx4));
assign Jeswx4 = (Qeswx4 & Xeswx4);
assign Xeswx4 = (~(Ohwvx4 & Mc9vx4));
assign Qeswx4 = (Efswx4 & Qpwvx4);
assign Qpwvx4 = (~(Mljwx4 & Ukpvx4));
assign Mljwx4 = (~(Zjwvx4 | Lcpvx4));
assign Efswx4 = (~(Nzgwx4 & Ukpvx4));
assign Nzgwx4 = (~(Zjwvx4 | Qfsvx4));
assign Zjwvx4 = (!V1yvx4);
assign V1yvx4 = (~(Iufwx4 | Kg9vx4));
assign Ceswx4 = (Z3yvx4 & Lfswx4);
assign Lfswx4 = (N4yvx4 | Mj8vx4);
assign Z3yvx4 = (Sfswx4 & Gkwvx4);
assign Gkwvx4 = (~(Pswvx4 & C2yvx4));
assign Pswvx4 = (~(Icyvx4 | Lcpvx4));
assign Sfswx4 = (~(Ohwvx4 & Epxvx4));
assign Odswx4 = (~(K79vx4 & Qslwx4));
assign Qslwx4 = (~(P7wvx4 & Zfswx4));
assign Zfswx4 = (~(Ukpvx4 & Pyxvx4));
assign Ukpvx4 = (Sh9vx4 & O4ovx4);
assign Pfhvx4 = (K6yvx4 ? Ggswx4 : Nt8vx4);
assign Ggswx4 = (~(Ngswx4 & Ugswx4));
assign Ugswx4 = (Bhswx4 & Ihswx4);
assign Ihswx4 = (Icyvx4 | J8svx4);
assign Bhswx4 = (Phswx4 & Whswx4);
assign Whswx4 = (~(H8yvx4 & I29vx4));
assign Phswx4 = (~(D69vx4 & Zayvx4));
assign Zayvx4 = (~(Iufwx4 & Diswx4));
assign Diswx4 = (Yj6wx4 | Fdsvx4);
assign Yj6wx4 = (!Ahwvx4);
assign Iufwx4 = (!Csewx4);
assign Ngswx4 = (Kiswx4 & G2lwx4);
assign Kiswx4 = (Riswx4 & Yiswx4);
assign Yiswx4 = (~(C9yvx4 & Layvx4));
assign Riswx4 = (~(Wv9vx4 & Pcyvx4));
assign Ifhvx4 = (K6yvx4 ? Fjswx4 : Vu8vx4);
assign K6yvx4 = (Mjswx4 & hready_i);
assign Mjswx4 = (~(Tjswx4 & Akswx4));
assign Akswx4 = (Hkswx4 & Okswx4);
assign Okswx4 = (Vkswx4 & Clswx4);
assign Clswx4 = (~(Jlswx4 & Ipkwx4));
assign Ipkwx4 = (Qlswx4 & Pyxvx4);
assign Pyxvx4 = (!Icyvx4);
assign Icyvx4 = (~(Xhxvx4 & Cf9vx4));
assign Qlswx4 = (~(Mj8vx4 | Aj9vx4));
assign Jlswx4 = (Xlswx4 & M1xvx4);
assign M1xvx4 = (!Ho8vx4);
assign Xlswx4 = (Sh9vx4 | U1fwx4);
assign U1fwx4 = (~(Qfsvx4 | Mc9vx4));
assign Vkswx4 = (Fhgwx4 & Tuwvx4);
assign Tuwvx4 = (~(Emswx4 & Lmswx4));
assign Lmswx4 = (~(Us2wx4 | Vdgvx4));
assign Emswx4 = (~(Ujxvx4 | Pxyvx4));
assign Fhgwx4 = (~(Zzfwx4 & Mcgvx4));
assign Hkswx4 = (Smswx4 & Zmswx4);
assign Zmswx4 = (~(D13wx4 & Gnswx4));
assign Gnswx4 = (W9fwx4 | Mj8vx4);
assign W9fwx4 = (!Rexvx4);
assign D13wx4 = (~(Hq1wx4 | Pxyvx4));
assign Smswx4 = (Nnswx4 & Unswx4);
assign Unswx4 = (~(Xlewx4 & Pkxvx4));
assign Xlewx4 = (~(Bl3wx4 | Mcgvx4));
assign Nnswx4 = (~(Ilpvx4 & Boswx4));
assign Boswx4 = (Ibdwx4 | Pa7wx4);
assign Pa7wx4 = (~(S87wx4 | U0ovx4));
assign Ilpvx4 = (Rngwx4 & Izwvx4);
assign Tjswx4 = (Ioswx4 & Poswx4);
assign Poswx4 = (Woswx4 & Dpswx4);
assign Dpswx4 = (X8kwx4 | Gwrvx4);
assign Gwrvx4 = (!P39vx4);
assign X8kwx4 = (~(Kpswx4 & Srgwx4));
assign Srgwx4 = (Rpswx4 & Ypswx4);
assign Ypswx4 = (~(Sh9vx4 | Mcgvx4));
assign Rpswx4 = (Howvx4 & K8hwx4);
assign Kpswx4 = (~(U4yvx4 | U9gvx4));
assign Woswx4 = (Fqswx4 & Mqswx4);
assign Mqswx4 = (~(Tqswx4 & O4ovx4));
assign Tqswx4 = (~(Arswx4 & Hrswx4));
assign Hrswx4 = (~(Orswx4 & C9yvx4));
assign Orswx4 = (~(Oedwx4 | Z6gvx4));
assign Arswx4 = (~(L5wvx4 & Sjwvx4));
assign Sjwvx4 = (Mgwvx4 & Sh9vx4);
assign L5wvx4 = (!X5gwx4);
assign X5gwx4 = (~(Xhxvx4 & Qfsvx4));
assign Xhxvx4 = (Cn8vx4 & Dfpvx4);
assign Fqswx4 = (~(Vrswx4 & Qfsvx4));
assign Qfsvx4 = (!Ud9vx4);
assign Vrswx4 = (~(Csswx4 & Jsswx4));
assign Jsswx4 = (~(Qsswx4 & Xsswx4));
assign Xsswx4 = (Etswx4 & Ejpvx4);
assign Ejpvx4 = (Y99vx4 & Cf9vx4);
assign Etswx4 = (~(Lqwvx4 | D69vx4));
assign Lqwvx4 = (!Dj6wx4);
assign Dj6wx4 = (~(Uasvx4 | Mc9vx4));
assign Qsswx4 = (~(J16wx4 | P7wvx4));
assign P7wvx4 = (~(Ltswx4 & Qsewx4));
assign Qsewx4 = (~(Dfpvx4 | Xmsvx4));
assign Ltswx4 = (Wvewx4 & O4ovx4);
assign Wvewx4 = (~(Lcpvx4 | Izwvx4));
assign J16wx4 = (!M4fwx4);
assign M4fwx4 = (~(Y5svx4 | K79vx4));
assign Y5svx4 = (!R89vx4);
assign Csswx4 = (~(Stswx4 & Ztswx4));
assign Ztswx4 = (~(Epxvx4 | Abgwx4));
assign Abgwx4 = (!G27wx4);
assign G27wx4 = (~(Uasvx4 | Fdsvx4));
assign Uasvx4 = (!Fb9vx4);
assign Epxvx4 = (!Jjgwx4);
assign Jjgwx4 = (~(Lcpvx4 | Bisvx4));
assign Stswx4 = (O3hwx4 & Ohwvx4);
assign Ohwvx4 = (Ahwvx4 & C2yvx4);
assign O3hwx4 = (Nywvx4 & J8svx4);
assign J8svx4 = (!Y99vx4);
assign Nywvx4 = (Zn6wx4 & D69vx4);
assign Ioswx4 = (I2mwx4 & Guswx4);
assign Guswx4 = (~(T1xvx4 & Ncqvx4));
assign I2mwx4 = (Lbiwx4 & Nuswx4);
assign Nuswx4 = (~(G0ovx4 & Clewx4));
assign G0ovx4 = (Ucqvx4 & Z6gvx4);
assign Fjswx4 = (~(Uuswx4 & Bvswx4));
assign Bvswx4 = (Ivswx4 & Pvswx4);
assign Pvswx4 = (~(H8yvx4 & P39vx4));
assign H8yvx4 = (Ahwvx4 & Fdsvx4);
assign Fdsvx4 = (!Mc9vx4);
assign Ivswx4 = (Wvswx4 & Dwswx4);
assign Dwswx4 = (~(Kwswx4 & Mc9vx4));
assign Kwswx4 = (K79vx4 & Rwswx4);
assign Rwswx4 = (Ahwvx4 | Csewx4);
assign Csewx4 = (~(Izwvx4 | Cf9vx4));
assign Ahwvx4 = (~(Dfpvx4 | Izwvx4));
assign Dfpvx4 = (!Kg9vx4);
assign Wvswx4 = (~(C9yvx4 & Ywswx4));
assign Ywswx4 = (~(Qmkwx4 & Fxswx4));
assign Fxswx4 = (~(Mxswx4 & Layvx4));
assign Mxswx4 = (~(Zrvvx4 | X0lwx4));
assign Qmkwx4 = (!Emewx4);
assign Emewx4 = (~(Q0lwx4 | Ks9vx4));
assign Uuswx4 = (G2lwx4 & Txswx4);
assign Txswx4 = (~(Bx9vx4 & Pcyvx4));
assign G2lwx4 = (Ayswx4 & Nbyvx4);
assign Nbyvx4 = (H2xvx4 & Vp2wx4);
assign Vp2wx4 = (~(Kzxvx4 & Dbgvx4));
assign H2xvx4 = (Pxyvx4 | B1ovx4);
assign Ayswx4 = (~(Zzfwx4 | Howvx4));
assign Bfhvx4 = (~(Hyswx4 & Oyswx4));
assign Oyswx4 = (Vyswx4 & Czswx4);
assign Czswx4 = (~(Xdfwx4 & Dmh2z4[9]));
assign Vyswx4 = (Jzswx4 & Lefwx4);
assign Jzswx4 = (Sefwx4 | Vq1wx4);
assign Vq1wx4 = (Qzswx4 & Xzswx4);
assign Xzswx4 = (E0twx4 & L0twx4);
assign L0twx4 = (~(Sknwx4 & Khfwx4));
assign Khfwx4 = (~(S0twx4 & Z0twx4));
assign Z0twx4 = (G1twx4 & N1twx4);
assign N1twx4 = (U1twx4 & B2twx4);
assign B2twx4 = (~(F9owx4 & L0i2z4[9]));
assign U1twx4 = (Ecowx4 & I2twx4);
assign G1twx4 = (P2twx4 & W2twx4);
assign W2twx4 = (~(M9owx4 & T1i2z4[9]));
assign P2twx4 = (~(Bzowx4 & Yxdwx4));
assign S0twx4 = (D3twx4 & K3twx4);
assign K3twx4 = (R3twx4 & Y3twx4);
assign Y3twx4 = (~(Fuowx4 & Zndwx4));
assign R3twx4 = (~(hrdata_i[9] & B7owx4));
assign D3twx4 = (F4twx4 & M4twx4);
assign M4twx4 = (~(Irh2z4[9] & I7owx4));
assign F4twx4 = (~(Czh2z4[9] & G6owx4));
assign E0twx4 = (T4twx4 & Glnwx4);
assign T4twx4 = (~(Pmnwx4 & Rhfwx4));
assign Rhfwx4 = (~(A5twx4 & H5twx4));
assign H5twx4 = (O5twx4 & V5twx4);
assign V5twx4 = (~(Bzowx4 & Fkdwx4));
assign O5twx4 = (C6twx4 & J6twx4);
assign J6twx4 = (~(H3owx4 & Q6twx4));
assign Q6twx4 = (~(X6twx4 & E7twx4));
assign E7twx4 = (L7twx4 & S7twx4);
assign S7twx4 = (~(S0hvx4 & A6tvx4));
assign A6tvx4 = (!A5uvx4);
assign A5uvx4 = (~(Z7twx4 & G8twx4));
assign Z7twx4 = (~(Z7hvx4 | L9hvx4));
assign L7twx4 = (~(T1i2z4[1] & Ts5wx4));
assign X6twx4 = (N8twx4 & U8twx4);
assign U8twx4 = (~(B2uvx4 & Eg8vx4));
assign N8twx4 = (~(M5tvx4 & L0i2z4[1]));
assign C6twx4 = (~(Fuowx4 & Jmdwx4));
assign A5twx4 = (B9twx4 & I9twx4);
assign I9twx4 = (~(Czh2z4[1] & G6owx4));
assign B9twx4 = (P9twx4 & W9twx4);
assign W9twx4 = (~(hrdata_i[1] & B7owx4));
assign P9twx4 = (~(Irh2z4[1] & I7owx4));
assign Qzswx4 = (Datwx4 & Katwx4);
assign Katwx4 = (~(Nlnwx4 & Bgfwx4));
assign Bgfwx4 = (~(Ratwx4 & Yatwx4));
assign Yatwx4 = (Fbtwx4 & Mbtwx4);
assign Mbtwx4 = (~(hrdata_i[17] & B7owx4));
assign Fbtwx4 = (Tbtwx4 & Actwx4);
assign Actwx4 = (~(Bzowx4 & Mrdwx4));
assign Tbtwx4 = (~(Fuowx4 & Jtdwx4));
assign Ratwx4 = (Hctwx4 & Octwx4);
assign Octwx4 = (~(Irh2z4[17] & I7owx4));
assign Hctwx4 = (~(Czh2z4[17] & G6owx4));
assign Datwx4 = (~(Imnwx4 & Pgfwx4));
assign Pgfwx4 = (~(Vctwx4 & Cdtwx4));
assign Cdtwx4 = (Jdtwx4 & T2owx4);
assign Jdtwx4 = (M7qwx4 | Qdtwx4);
assign Vctwx4 = (Xdtwx4 & Eetwx4);
assign Eetwx4 = (~(M5ewx4 & L5owx4));
assign M5ewx4 = (Letwx4 & Qdtwx4);
assign Qdtwx4 = (Setwx4 | V8qwx4);
assign Setwx4 = (Zetwx4 ? Udowx4 : C9qwx4);
assign Letwx4 = (Yw7wx4 ? Gftwx4 : Gvdwx4);
assign Xdtwx4 = (~(hrdata_i[25] & B7owx4));
assign Hyswx4 = (Nftwx4 & Uftwx4);
assign Uftwx4 = (~(Roh2z4[8] & Mifwx4));
assign Nftwx4 = (~(vis_pc_o[8] & Qaiwx4));
assign Uehvx4 = (~(Bgtwx4 & Igtwx4));
assign Igtwx4 = (Pgtwx4 & Wgtwx4);
assign Wgtwx4 = (~(Xdfwx4 & Dmh2z4[11]));
assign Pgtwx4 = (Dhtwx4 & Lefwx4);
assign Dhtwx4 = (Sefwx4 | Ll1wx4);
assign Ll1wx4 = (Khtwx4 & Rhtwx4);
assign Rhtwx4 = (Yhtwx4 & Fitwx4);
assign Fitwx4 = (~(Sknwx4 & Whlwx4));
assign Whlwx4 = (~(Mitwx4 & Titwx4));
assign Titwx4 = (Ajtwx4 & Hjtwx4);
assign Hjtwx4 = (Ojtwx4 & Vjtwx4);
assign Vjtwx4 = (~(F9owx4 & L0i2z4[11]));
assign Ojtwx4 = (~(M9owx4 & T1i2z4[11]));
assign Ajtwx4 = (Cktwx4 & Jktwx4);
assign Jktwx4 = (~(Fuowx4 & Vzdwx4));
assign Cktwx4 = (~(Bzowx4 & X0ewx4));
assign Mitwx4 = (Qktwx4 & Xktwx4);
assign Xktwx4 = (~(Czh2z4[11] & G6owx4));
assign Qktwx4 = (Eltwx4 & Lltwx4);
assign Lltwx4 = (~(hrdata_i[11] & B7owx4));
assign Eltwx4 = (~(Irh2z4[11] & I7owx4));
assign Yhtwx4 = (Sltwx4 & Glnwx4);
assign Sltwx4 = (~(Pmnwx4 & Ihlwx4));
assign Ihlwx4 = (~(Zltwx4 & Gmtwx4));
assign Gmtwx4 = (Nmtwx4 & Umtwx4);
assign Umtwx4 = (Bntwx4 & I2twx4);
assign I2twx4 = (~(Intwx4 & Pntwx4));
assign Pntwx4 = (Wntwx4 & Z7hvx4);
assign Wntwx4 = (~(B5hvx4 | L9hvx4));
assign Intwx4 = (H3owx4 & Dotwx4);
assign Bntwx4 = (~(F9owx4 & L0i2z4[3]));
assign Nmtwx4 = (Kotwx4 & Rotwx4);
assign Rotwx4 = (~(M9owx4 & T1i2z4[3]));
assign Kotwx4 = (~(Bzowx4 & Nodwx4));
assign Zltwx4 = (Yotwx4 & Fptwx4);
assign Fptwx4 = (Mptwx4 & Tptwx4);
assign Tptwx4 = (~(Fuowx4 & Rw7wx4));
assign Mptwx4 = (~(hrdata_i[3] & B7owx4));
assign Yotwx4 = (Aqtwx4 & Hqtwx4);
assign Hqtwx4 = (~(Irh2z4[3] & I7owx4));
assign Aqtwx4 = (~(Czh2z4[3] & G6owx4));
assign Khtwx4 = (Oqtwx4 & Vqtwx4);
assign Vqtwx4 = (~(Nlnwx4 & Rilwx4));
assign Rilwx4 = (~(Crtwx4 & Jrtwx4));
assign Jrtwx4 = (Qrtwx4 & Xrtwx4);
assign Xrtwx4 = (~(Fuowx4 & Qtdwx4));
assign Qrtwx4 = (Estwx4 & Ecowx4);
assign Ecowx4 = (X3pwx4 | Lstwx4);
assign Estwx4 = (~(Bzowx4 & Uvdwx4));
assign Crtwx4 = (Sstwx4 & Zstwx4);
assign Zstwx4 = (~(Czh2z4[19] & G6owx4));
assign Sstwx4 = (Gttwx4 & Nttwx4);
assign Nttwx4 = (~(hrdata_i[19] & B7owx4));
assign Gttwx4 = (~(Irh2z4[19] & I7owx4));
assign Oqtwx4 = (~(Imnwx4 & Mjlwx4));
assign Mjlwx4 = (~(Uttwx4 & Butwx4));
assign Butwx4 = (Iutwx4 & T2owx4);
assign Iutwx4 = (~(H6ewx4 & Putwx4));
assign Putwx4 = (Fuowx4 | Wutwx4);
assign Wutwx4 = (L5owx4 & Kw7wx4);
assign H6ewx4 = (Dvtwx4 & Kvtwx4);
assign Dvtwx4 = (~(Rvtwx4 & Yvtwx4));
assign Rvtwx4 = (Oldwx4 & Fwtwx4);
assign Uttwx4 = (Mwtwx4 & Twtwx4);
assign Twtwx4 = (Kvtwx4 | M7qwx4);
assign Kvtwx4 = (Axtwx4 | V8qwx4);
assign V8qwx4 = (~(Mcgvx4 & Weowx4));
assign Axtwx4 = (A1qwx4 ? C9qwx4 : Udowx4);
assign Mwtwx4 = (~(hrdata_i[27] & B7owx4));
assign Bgtwx4 = (Hxtwx4 & Oxtwx4);
assign Oxtwx4 = (~(Roh2z4[10] & Mifwx4));
assign Hxtwx4 = (~(vis_pc_o[10] & Qaiwx4));
assign Nehvx4 = (~(Vxtwx4 & Cytwx4));
assign Cytwx4 = (Jytwx4 & Qytwx4);
assign Qytwx4 = (~(Xdfwx4 & Dmh2z4[13]));
assign Jytwx4 = (Xytwx4 & Lefwx4);
assign Xytwx4 = (Sefwx4 | Mb1wx4);
assign Mb1wx4 = (Eztwx4 & Lztwx4);
assign Lztwx4 = (Sztwx4 & Zztwx4);
assign Zztwx4 = (~(Sknwx4 & Twmwx4));
assign Sztwx4 = (G0uwx4 & Glnwx4);
assign G0uwx4 = (~(Nlnwx4 & Jymwx4));
assign Eztwx4 = (N0uwx4 & U0uwx4);
assign U0uwx4 = (~(Imnwx4 & Hxmwx4));
assign N0uwx4 = (~(Pmnwx4 & Cymwx4));
assign Vxtwx4 = (B1uwx4 & I1uwx4);
assign I1uwx4 = (~(Roh2z4[12] & Mifwx4));
assign B1uwx4 = (~(vis_pc_o[12] & Qaiwx4));
assign Gehvx4 = (~(P1uwx4 & W1uwx4));
assign W1uwx4 = (D2uwx4 & K2uwx4);
assign K2uwx4 = (~(Roh2z4[20] & Mifwx4));
assign D2uwx4 = (R2uwx4 & Y2uwx4);
assign Y2uwx4 = (Sefwx4 | Qe0wx4);
assign Qe0wx4 = (F3uwx4 & M3uwx4);
assign M3uwx4 = (T3uwx4 & A4uwx4);
assign A4uwx4 = (~(Jymwx4 & Yilwx4));
assign Jymwx4 = (~(H4uwx4 & O4uwx4));
assign O4uwx4 = (V4uwx4 & C5uwx4);
assign C5uwx4 = (~(hrdata_i[21] & B7owx4));
assign V4uwx4 = (J5uwx4 & Q5uwx4);
assign Q5uwx4 = (~(Bzowx4 & Gvdwx4));
assign Gvdwx4 = (~(X5uwx4 & E6uwx4));
assign E6uwx4 = (L6uwx4 & S6uwx4);
assign S6uwx4 = (~(O1qwx4 & Kdqwx4));
assign L6uwx4 = (~(Yzpwx4 & Z6uwx4));
assign X5uwx4 = (G7uwx4 & N7uwx4);
assign N7uwx4 = (A1qwx4 | U7uwx4);
assign G7uwx4 = (~(Kzpwx4 & Meqwx4));
assign J5uwx4 = (~(Fuowx4 & Mrdwx4));
assign Mrdwx4 = (~(B8uwx4 & I8uwx4));
assign I8uwx4 = (P8uwx4 & W8uwx4);
assign W8uwx4 = (~(O1qwx4 & N4qwx4));
assign P8uwx4 = (A1qwx4 | D9uwx4);
assign B8uwx4 = (K9uwx4 & R9uwx4);
assign R9uwx4 = (~(Yzpwx4 & Y9uwx4));
assign K9uwx4 = (~(Kzpwx4 & L3qwx4));
assign H4uwx4 = (Fauwx4 & Mauwx4);
assign Mauwx4 = (~(Irh2z4[21] & I7owx4));
assign Fauwx4 = (~(Czh2z4[21] & G6owx4));
assign T3uwx4 = (~(Phlwx4 & Twmwx4));
assign Twmwx4 = (~(Tauwx4 & Abuwx4));
assign Abuwx4 = (Hbuwx4 & Obuwx4);
assign Obuwx4 = (~(Bzowx4 & Jtdwx4));
assign Jtdwx4 = (~(Vbuwx4 & Ccuwx4));
assign Ccuwx4 = (Jcuwx4 & Qcuwx4);
assign Qcuwx4 = (~(O1qwx4 & F0qwx4));
assign Jcuwx4 = (A1qwx4 | Xcuwx4);
assign Vbuwx4 = (Eduwx4 & Lduwx4);
assign Lduwx4 = (~(Yzpwx4 & Sduwx4));
assign Eduwx4 = (~(Kzpwx4 & V1qwx4));
assign Hbuwx4 = (Zduwx4 & Geuwx4);
assign Geuwx4 = (~(H3owx4 & Neuwx4));
assign Neuwx4 = (~(Ueuwx4 & Bfuwx4));
assign Bfuwx4 = (~(M5tvx4 & L0i2z4[13]));
assign Ueuwx4 = (Ifuwx4 & Pfuwx4);
assign Pfuwx4 = (Wfuwx4 | Kzqvx4);
assign Kzqvx4 = (Dguwx4 & Kguwx4);
assign Kguwx4 = (~(Rguwx4 & Yguwx4));
assign Rguwx4 = (~(Fhuwx4 & Mhuwx4));
assign Mhuwx4 = (I6pwx4 ? Aiuwx4 : Thuwx4);
assign Aiuwx4 = (~(Hiuwx4 | Oiuwx4));
assign Oiuwx4 = (~(B6pwx4 | Viuwx4));
assign Thuwx4 = (U5pwx4 ? Jjuwx4 : Cjuwx4);
assign Fhuwx4 = (Qjuwx4 & G5pwx4);
assign Ifuwx4 = (~(T1i2z4[13] & Ts5wx4));
assign Zduwx4 = (~(Fuowx4 & Yxdwx4));
assign Yxdwx4 = (~(Xjuwx4 & Ekuwx4));
assign Ekuwx4 = (Lkuwx4 & Skuwx4);
assign Skuwx4 = (~(O1qwx4 & Omqwx4));
assign Lkuwx4 = (A1qwx4 | Zkuwx4);
assign Xjuwx4 = (Gluwx4 & Nluwx4);
assign Nluwx4 = (~(Yzpwx4 & Uluwx4));
assign Gluwx4 = (~(Kzpwx4 & Mlqwx4));
assign Tauwx4 = (Bmuwx4 & Imuwx4);
assign Imuwx4 = (~(Czh2z4[13] & G6owx4));
assign Bmuwx4 = (Pmuwx4 & Wmuwx4);
assign Wmuwx4 = (~(hrdata_i[13] & B7owx4));
assign Pmuwx4 = (~(Irh2z4[13] & I7owx4));
assign F3uwx4 = (Dnuwx4 & Knuwx4);
assign Knuwx4 = (~(Fjlwx4 & Hxmwx4));
assign Hxmwx4 = (~(Rnuwx4 & Ynuwx4));
assign Ynuwx4 = (Fouwx4 & T2owx4);
assign Fouwx4 = (Mouwx4 | M7qwx4);
assign M7qwx4 = (~(U2ewx4 & L5owx4));
assign Rnuwx4 = (Touwx4 & Apuwx4);
assign Apuwx4 = (~(F5ewx4 & L5owx4));
assign F5ewx4 = (Hpuwx4 & Mouwx4);
assign Mouwx4 = (~(Opuwx4 & Wdpwx4));
assign Opuwx4 = (Zetwx4 ? Weowx4 : Udowx4);
assign Zetwx4 = (Depwx4 | O1qwx4);
assign Depwx4 = (Yzpwx4 | Vpuwx4);
assign Hpuwx4 = (Oldwx4 ? Gftwx4 : Jmdwx4);
assign Gftwx4 = (~(Cquwx4 & Jquwx4));
assign Jquwx4 = (Qquwx4 & Xquwx4);
assign Xquwx4 = (~(O1qwx4 & Nbqwx4));
assign Qquwx4 = (A1qwx4 | Eruwx4);
assign Cquwx4 = (Lruwx4 & Sruwx4);
assign Sruwx4 = (~(Yzpwx4 & Zruwx4));
assign Lruwx4 = (~(Kzpwx4 & Laqwx4));
assign Jmdwx4 = (~(Gsuwx4 & Nsuwx4));
assign Nsuwx4 = (Usuwx4 & Btuwx4);
assign Btuwx4 = (~(O1qwx4 & Iqqwx4));
assign Usuwx4 = (~(Yzpwx4 & Ituwx4));
assign Gsuwx4 = (Ptuwx4 & Wtuwx4);
assign Wtuwx4 = (A1qwx4 | Duuwx4);
assign Ptuwx4 = (~(Kzpwx4 & Drqwx4));
assign Touwx4 = (~(hrdata_i[29] & B7owx4));
assign Dnuwx4 = (~(W6iwx4 & Cymwx4));
assign Cymwx4 = (~(Kuuwx4 & Ruuwx4));
assign Ruuwx4 = (Yuuwx4 & Fvuwx4);
assign Fvuwx4 = (Mvuwx4 & Tvuwx4);
assign Tvuwx4 = (~(F9owx4 & L0i2z4[5]));
assign F9owx4 = (H3owx4 & M5tvx4);
assign Mvuwx4 = (~(M9owx4 & T1i2z4[5]));
assign M9owx4 = (H3owx4 & Ts5wx4);
assign Yuuwx4 = (Awuwx4 & Hwuwx4);
assign Hwuwx4 = (~(Fuowx4 & Fkdwx4));
assign Fkdwx4 = (~(Owuwx4 & Vwuwx4));
assign Vwuwx4 = (Cxuwx4 & Jxuwx4);
assign Jxuwx4 = (~(O1qwx4 & Zvqwx4));
assign Cxuwx4 = (A1qwx4 | Qxuwx4);
assign Owuwx4 = (Xxuwx4 & Eyuwx4);
assign Eyuwx4 = (~(Yzpwx4 & Lyuwx4));
assign Xxuwx4 = (~(Kzpwx4 & Xuqwx4));
assign Awuwx4 = (~(Bzowx4 & Zndwx4));
assign Zndwx4 = (~(Syuwx4 & Zyuwx4));
assign Zyuwx4 = (Gzuwx4 & Nzuwx4);
assign Nzuwx4 = (~(O1qwx4 & Uiqwx4));
assign Gzuwx4 = (A1qwx4 | Pybwx4);
assign Syuwx4 = (Uzuwx4 & B0vwx4);
assign B0vwx4 = (~(Yzpwx4 & I0vwx4));
assign Uzuwx4 = (~(Kzpwx4 & Wjqwx4));
assign Kuuwx4 = (P0vwx4 & W0vwx4);
assign W0vwx4 = (~(Czh2z4[5] & G6owx4));
assign P0vwx4 = (D1vwx4 & K1vwx4);
assign K1vwx4 = (~(hrdata_i[5] & B7owx4));
assign D1vwx4 = (~(Irh2z4[5] & I7owx4));
assign R2uwx4 = (~(Xdfwx4 & Dmh2z4[21]));
assign P1uwx4 = (Tjlwx4 & R1vwx4);
assign R1vwx4 = (~(vis_pc_o[20] & Qaiwx4));
assign Zdhvx4 = (~(Y1vwx4 & F2vwx4));
assign F2vwx4 = (M2vwx4 & T2vwx4);
assign T2vwx4 = (~(Xdfwx4 & Dmh2z4[23]));
assign M2vwx4 = (A3vwx4 & Lefwx4);
assign A3vwx4 = (Sefwx4 | Oa3wx4);
assign Oa3wx4 = (H3vwx4 & O3vwx4);
assign O3vwx4 = (V3vwx4 & C4vwx4);
assign C4vwx4 = (~(W6iwx4 & G9lwx4));
assign V3vwx4 = (J4vwx4 & D31wx4);
assign J4vwx4 = (~(Yilwx4 & Walwx4));
assign H3vwx4 = (Q4vwx4 & X4vwx4);
assign X4vwx4 = (~(Fjlwx4 & Palwx4));
assign Q4vwx4 = (~(Phlwx4 & U9lwx4));
assign Y1vwx4 = (E5vwx4 & L5vwx4);
assign L5vwx4 = (~(Roh2z4[22] & Mifwx4));
assign E5vwx4 = (~(vis_pc_o[22] & Qaiwx4));
assign Sdhvx4 = (~(S5vwx4 & Z5vwx4));
assign Z5vwx4 = (G6vwx4 & N6vwx4);
assign N6vwx4 = (~(Xdfwx4 & Dmh2z4[15]));
assign G6vwx4 = (U6vwx4 & Lefwx4);
assign U6vwx4 = (Sefwx4 | U72wx4);
assign U72wx4 = (B7vwx4 & I7vwx4);
assign I7vwx4 = (P7vwx4 & W7vwx4);
assign W7vwx4 = (~(Sknwx4 & U9lwx4));
assign Sknwx4 = (~(Tanwx4 & D8vwx4));
assign D8vwx4 = (~(E6nwx4 & K8vwx4));
assign K8vwx4 = (~(K7xvx4 & R8vwx4));
assign R8vwx4 = (~(Y8vwx4 & N7nwx4));
assign Y8vwx4 = (~(O33wx4 & F9vwx4));
assign F9vwx4 = (H33wx4 | U9gvx4);
assign K7xvx4 = (!Wdqvx4);
assign Tanwx4 = (~(Yilwx4 | M9vwx4));
assign M9vwx4 = (T9vwx4 & E6nwx4);
assign T9vwx4 = (Ri7wx4 & Mcgvx4);
assign Ri7wx4 = (Nggvx4 & Dbgvx4);
assign P7vwx4 = (Aavwx4 & Glnwx4);
assign Glnwx4 = (~(B8nwx4 & Havwx4));
assign Havwx4 = (~(Oavwx4 & W8nwx4));
assign Oavwx4 = (R9nwx4 ? I3ewx4 : Vavwx4);
assign I3ewx4 = (~(Bwdwx4 & S1ewx4));
assign Bwdwx4 = (Fanwx4 & Qs7wx4);
assign Fanwx4 = (Bpdwx4 & Cbvwx4);
assign Vavwx4 = (Jbvwx4 & Qbvwx4);
assign Qbvwx4 = (~(Xbvwx4 & B1vvx4));
assign Xbvwx4 = (~(Izwvx4 | U9gvx4));
assign Jbvwx4 = (Y47wx4 | W5yvx4);
assign Aavwx4 = (~(Pmnwx4 & G9lwx4));
assign Pmnwx4 = (F8iwx4 | Ygnwx4);
assign Ygnwx4 = (Ecvwx4 & E6nwx4);
assign Ecvwx4 = (Wdxvx4 & Hw2wx4);
assign F8iwx4 = (~(Kgnwx4 & Lcvwx4));
assign B7vwx4 = (Scvwx4 & Zcvwx4);
assign Zcvwx4 = (~(Nlnwx4 & Walwx4));
assign Nlnwx4 = (~(Uenwx4 & Dgnwx4));
assign Dgnwx4 = (Cbvwx4 | E6nwx4);
assign Cbvwx4 = (Gdvwx4 | Y9nwx4);
assign Scvwx4 = (~(Imnwx4 & Palwx4));
assign Imnwx4 = (Ndvwx4 | S6nwx4);
assign S6nwx4 = (Udvwx4 & Bevwx4);
assign Bevwx4 = (~(Agqvx4 | B1ovx4));
assign Udvwx4 = (~(R9nwx4 | N7nwx4));
assign Ndvwx4 = (R9nwx4 ? Mq7wx4 : Ievwx4);
assign Ievwx4 = (~(O33wx4 | N7nwx4));
assign O33wx4 = (M3ovx4 | Dbgvx4);
assign S5vwx4 = (Pevwx4 & Wevwx4);
assign Wevwx4 = (~(Roh2z4[14] & Mifwx4));
assign Pevwx4 = (~(vis_pc_o[14] & Qaiwx4));
assign Ldhvx4 = (~(Dfvwx4 & Kfvwx4));
assign Kfvwx4 = (Rfvwx4 & Yfvwx4);
assign Yfvwx4 = (~(Roh2z4[19] & Mifwx4));
assign Mifwx4 = (~(S5pvx4 | Qaiwx4));
assign S5pvx4 = (M9pvx4 | Y8pvx4);
assign Rfvwx4 = (Fgvwx4 & Mgvwx4);
assign Mgvwx4 = (Sefwx4 | Tj0wx4);
assign Tj0wx4 = (Tgvwx4 & Ahvwx4);
assign Ahvwx4 = (Hhvwx4 & Ohvwx4);
assign Ohvwx4 = (~(Ntmwx4 & Yilwx4));
assign Yilwx4 = (~(S9rwx4 & Vhvwx4));
assign S9rwx4 = (~(E6nwx4 & Civwx4));
assign Civwx4 = (~(Cn8vx4 & Jivwx4));
assign Jivwx4 = (~(Tv2wx4 & Qivwx4));
assign Qivwx4 = (S4xvx4 | B1ovx4);
assign Ntmwx4 = (~(Xivwx4 & Ejvwx4));
assign Ejvwx4 = (Ljvwx4 & Sjvwx4);
assign Sjvwx4 = (~(hrdata_i[20] & B7owx4));
assign Ljvwx4 = (Zjvwx4 & Gkvwx4);
assign Gkvwx4 = (~(Fuowx4 & Xtdwx4));
assign Xtdwx4 = (~(Nkvwx4 & Ukvwx4));
assign Ukvwx4 = (Blvwx4 & Ilvwx4);
assign Ilvwx4 = (~(O1qwx4 & Y9uwx4));
assign Blvwx4 = (~(Kzpwx4 & N4qwx4));
assign Nkvwx4 = (Plvwx4 & Wlvwx4);
assign Wlvwx4 = (~(Yzpwx4 & Rzpwx4));
assign Plvwx4 = (A1qwx4 | Dmvwx4);
assign Zjvwx4 = (~(Bzowx4 & Nvdwx4));
assign Nvdwx4 = (~(Kmvwx4 & Rmvwx4));
assign Rmvwx4 = (Ymvwx4 & Fnvwx4);
assign Fnvwx4 = (~(O1qwx4 & Z6uwx4));
assign Ymvwx4 = (A1qwx4 | Mnvwx4);
assign Kmvwx4 = (Tnvwx4 & Aovwx4);
assign Aovwx4 = (~(Yzpwx4 & E3qwx4));
assign Tnvwx4 = (~(Kzpwx4 & Kdqwx4));
assign Xivwx4 = (Hovwx4 & Oovwx4);
assign Oovwx4 = (~(Irh2z4[20] & I7owx4));
assign Hovwx4 = (~(Czh2z4[20] & G6owx4));
assign Hhvwx4 = (~(Phlwx4 & Xrmwx4));
assign Xrmwx4 = (~(Vovwx4 & Cpvwx4));
assign Cpvwx4 = (Jpvwx4 & Qpvwx4);
assign Qpvwx4 = (~(Bzowx4 & E1ewx4));
assign E1ewx4 = (~(Xpvwx4 & Eqvwx4));
assign Eqvwx4 = (Lqvwx4 & Sqvwx4);
assign Sqvwx4 = (~(O1qwx4 & Sduwx4));
assign Lqvwx4 = (~(Kzpwx4 & F0qwx4));
assign Xpvwx4 = (Zqvwx4 & Grvwx4);
assign Grvwx4 = (~(Yzpwx4 & Flqwx4));
assign Zqvwx4 = (A1qwx4 | Nrvwx4);
assign Jpvwx4 = (Urvwx4 & Bsvwx4);
assign Bsvwx4 = (~(H3owx4 & Isvwx4));
assign Isvwx4 = (~(Psvwx4 & Wsvwx4));
assign Wsvwx4 = (~(M5tvx4 & L0i2z4[12]));
assign Psvwx4 = (Dtvwx4 & Ktvwx4);
assign Ktvwx4 = (Ewqvx4 | Wfuwx4);
assign Ewqvx4 = (!Kkrvx4);
assign Kkrvx4 = (Rtvwx4 & Sw4wx4);
assign Rtvwx4 = (~(Ytvwx4 & Fuvwx4));
assign Fuvwx4 = (Muvwx4 | Tuvwx4);
assign Tuvwx4 = (!Yguwx4);
assign Muvwx4 = (G5pwx4 ? Hvvwx4 : Avvwx4);
assign Hvvwx4 = (Qjuwx4 & Ovvwx4);
assign Ovvwx4 = (I6pwx4 ? Cwvwx4 : Vvvwx4);
assign Cwvwx4 = (Jwvwx4 & Qwvwx4);
assign Qwvwx4 = (~(Hiuwx4 & Xwvwx4));
assign Jwvwx4 = (B6pwx4 ? Lxvwx4 : Exvwx4);
assign Lxvwx4 = (Sxvwx4 | Zxvwx4);
assign Exvwx4 = (Viuwx4 ? Nyvwx4 : Gyvwx4);
assign Vvvwx4 = (U5pwx4 ? Bzvwx4 : Uyvwx4);
assign Bzvwx4 = (!Izvwx4);
assign Izvwx4 = (Jjuwx4 ? Wzvwx4 : Pzvwx4);
assign Uyvwx4 = (Cjuwx4 ? K0wwx4 : D0wwx4);
assign Dtvwx4 = (~(T1i2z4[12] & Ts5wx4));
assign Urvwx4 = (~(Fuowx4 & C0ewx4));
assign C0ewx4 = (~(R0wwx4 & Y0wwx4));
assign Y0wwx4 = (F1wwx4 & M1wwx4);
assign M1wwx4 = (~(O1qwx4 & Uluwx4));
assign F1wwx4 = (~(Kzpwx4 & Omqwx4));
assign R0wwx4 = (T1wwx4 & A2wwx4);
assign A2wwx4 = (~(Yzpwx4 & Niqwx4));
assign T1wwx4 = (A1qwx4 | H2wwx4);
assign Vovwx4 = (O2wwx4 & V2wwx4);
assign V2wwx4 = (~(Czh2z4[12] & G6owx4));
assign O2wwx4 = (C3wwx4 & J3wwx4);
assign J3wwx4 = (~(hrdata_i[12] & B7owx4));
assign C3wwx4 = (~(Irh2z4[12] & I7owx4));
assign Phlwx4 = (~(Uenwx4 & Lcvwx4));
assign Uenwx4 = (R9nwx4 | M93wx4);
assign R9nwx4 = (!E6nwx4);
assign Tgvwx4 = (Q3wwx4 & X3wwx4);
assign X3wwx4 = (~(Fjlwx4 & Lsmwx4));
assign Lsmwx4 = (~(E4wwx4 & L4wwx4));
assign L4wwx4 = (S4wwx4 & T2owx4);
assign T2owx4 = (~(Z4wwx4 & H3owx4));
assign S4wwx4 = (~(C4owx4 & Qsgvx4));
assign C4owx4 = (H3owx4 & Gc4wx4);
assign E4wwx4 = (G5wwx4 & N5wwx4);
assign N5wwx4 = (Lcowx4 | X7ewx4);
assign X7ewx4 = (U5wwx4 & B6wwx4);
assign B6wwx4 = (~(I6wwx4 & U2ewx4));
assign I6wwx4 = (Wdpwx4 & Weowx4);
assign U5wwx4 = (~(P6wwx4 & W6wwx4));
assign W6wwx4 = (~(Wdpwx4 & Weowx4));
assign P6wwx4 = (Oldwx4 ? Beowx4 : Jiowx4);
assign Beowx4 = (~(D7wwx4 & K7wwx4));
assign K7wwx4 = (R7wwx4 & Y7wwx4);
assign Y7wwx4 = (~(O1qwx4 & Zruwx4));
assign R7wwx4 = (A1qwx4 | F8wwx4);
assign D7wwx4 = (M8wwx4 & T8wwx4);
assign T8wwx4 = (~(Yzpwx4 & Ddqwx4));
assign M8wwx4 = (~(Kzpwx4 & Nbqwx4));
assign Jiowx4 = (~(A9wwx4 & H9wwx4));
assign H9wwx4 = (O9wwx4 & V9wwx4);
assign V9wwx4 = (~(O1qwx4 & Ituwx4));
assign O9wwx4 = (A1qwx4 | Cawwx4);
assign A9wwx4 = (Jawwx4 & Qawwx4);
assign Qawwx4 = (~(Yzpwx4 & Ubqwx4));
assign Jawwx4 = (~(Kzpwx4 & Iqqwx4));
assign G5wwx4 = (~(hrdata_i[28] & B7owx4));
assign Fjlwx4 = (~(Kgnwx4 & C8rwx4));
assign Kgnwx4 = (~(E6nwx4 & Jp3wx4));
assign Q3wwx4 = (~(W6iwx4 & Gtmwx4));
assign Gtmwx4 = (~(Xawwx4 & Ebwwx4));
assign Ebwwx4 = (Lbwwx4 & Sbwwx4);
assign Sbwwx4 = (~(Fuowx4 & Qmdwx4));
assign Qmdwx4 = (~(Zbwwx4 & Gcwwx4));
assign Gcwwx4 = (Ncwwx4 & Ucwwx4);
assign Ucwwx4 = (~(O1qwx4 & Lyuwx4));
assign Ncwwx4 = (A1qwx4 | Bdwwx4);
assign Zbwwx4 = (Idwwx4 & Pdwwx4);
assign Pdwwx4 = (~(Yzpwx4 & Bqqwx4));
assign Idwwx4 = (~(Kzpwx4 & Zvqwx4));
assign Fuowx4 = (~(Lcowx4 | Yw7wx4));
assign Lbwwx4 = (Wdwwx4 & Dewwx4);
assign Dewwx4 = (~(H3owx4 & Kewwx4));
assign Kewwx4 = (~(Rewwx4 & Yewwx4));
assign Yewwx4 = (~(M5tvx4 & L0i2z4[4]));
assign Rewwx4 = (Ffwwx4 & Mfwwx4);
assign Mfwwx4 = (~(T1i2z4[4] & Ts5wx4));
assign Ffwwx4 = (~(Vogvx4 & B2uvx4));
assign B2uvx4 = (Vssvx4 & Z7hvx4);
assign Wdwwx4 = (~(hrdata_i[4] & B7owx4));
assign Xawwx4 = (Tfwwx4 & Agwwx4);
assign Agwwx4 = (~(Czh2z4[4] & G6owx4));
assign Tfwwx4 = (Hgwwx4 & Ogwwx4);
assign Ogwwx4 = (~(Irh2z4[4] & I7owx4));
assign Hgwwx4 = (~(Bzowx4 & Godwx4));
assign Godwx4 = (~(Vgwwx4 & Chwwx4));
assign Chwwx4 = (Jhwwx4 & Qhwwx4);
assign Qhwwx4 = (~(O1qwx4 & I0vwx4));
assign Jhwwx4 = (~(Kzpwx4 & Uiqwx4));
assign Vgwwx4 = (Xhwwx4 & Eiwwx4);
assign Eiwwx4 = (~(Yzpwx4 & Quqwx4));
assign Xhwwx4 = (A1qwx4 | Lr9wx4);
assign Bzowx4 = (L5owx4 & Yw7wx4);
assign Fgvwx4 = (~(Xdfwx4 & Dmh2z4[20]));
assign Xdfwx4 = (G6pvx4 & M9pvx4);
assign Dfvwx4 = (Tjlwx4 & Liwwx4);
assign Liwwx4 = (~(vis_pc_o[19] & Qaiwx4));
assign Tjlwx4 = (Lefwx4 & Siwwx4);
assign Siwwx4 = (D31wx4 | Sefwx4);
assign Sefwx4 = (!H4nwx4);
assign H4nwx4 = (G6pvx4 & Y8pvx4);
assign D31wx4 = (~(Ziwwx4 & Gjwwx4));
assign Gjwwx4 = (Njwwx4 & C8rwx4);
assign C8rwx4 = (Gdvwx4 | E6nwx4);
assign Gdvwx4 = (!Yp7wx4);
assign Yp7wx4 = (Ujwwx4 & Vy7wx4);
assign Ujwwx4 = (Cz7wx4 & Manwx4);
assign Njwwx4 = (~(Bkwwx4 | W6iwx4));
assign W6iwx4 = (Ikwwx4 & Mq7wx4);
assign Mq7wx4 = (!S1ewx4);
assign S1ewx4 = (~(Fx7wx4 & Manwx4));
assign Fx7wx4 = (~(Cz7wx4 | Vy7wx4));
assign Cz7wx4 = (!Pkwwx4);
assign Ikwwx4 = (~(Z1ewx4 | E6nwx4));
assign Bkwwx4 = (!Lcvwx4);
assign Lcvwx4 = (Qs7wx4 | E6nwx4);
assign Qs7wx4 = (~(Wkwwx4 & Ay7wx4));
assign Ay7wx4 = (~(Vy7wx4 | Pkwwx4));
assign Wkwwx4 = (Dp7wx4 & Manwx4);
assign Ziwwx4 = (Q8rwx4 & Vhvwx4);
assign Vhvwx4 = (Bpdwx4 | E6nwx4);
assign Bpdwx4 = (S8ewx4 | Y9nwx4);
assign Y9nwx4 = (~(F3ovx4 | Dlwwx4));
assign Dlwwx4 = (!Klwwx4);
assign S8ewx4 = (~(Dw7wx4 & Manwx4));
assign Manwx4 = (~(Mcgvx4 & Zm7wx4));
assign Zm7wx4 = (!Ok7wx4);
assign Ok7wx4 = (Rlwwx4 & Ylwwx4);
assign Ylwwx4 = (~(Fmwwx4 & Mmwwx4));
assign Mmwwx4 = (Tmwwx4 & U5bwx4);
assign U5bwx4 = (!Un9vx4);
assign Tmwwx4 = (~(Yo9vx4 | Z6gvx4));
assign Fmwwx4 = (Anwwx4 & Hnwwx4);
assign Anwwx4 = (Onwwx4 & Yryvx4);
assign Rlwwx4 = (Vnwwx4 & Gu7wx4);
assign Gu7wx4 = (~(Cowwx4 & Jowwx4));
assign Jowwx4 = (~(Qowwx4 & Xowwx4));
assign Vnwwx4 = (~(Cowwx4 & Epwwx4));
assign Epwwx4 = (~(Lpwwx4 & Spwwx4));
assign Lpwwx4 = (Zpwwx4 & Gqwwx4);
assign Q8rwx4 = (Nqwwx4 & B8nwx4);
assign B8nwx4 = (~(Uqwwx4 & Brwwx4));
assign Brwwx4 = (Irwwx4 & Prwwx4);
assign Prwwx4 = (~(Wrwwx4 & Wxcwx4));
assign Wrwwx4 = (~(Dswwx4 | U9gvx4));
assign Irwwx4 = (Kswwx4 & Js7wx4);
assign Js7wx4 = (!U2ewx4);
assign Kswwx4 = (~(Rswwx4 & Oe6wx4));
assign Oe6wx4 = (Whgvx4 & Nggvx4);
assign Rswwx4 = (Mcgvx4 & U9lwx4);
assign Uqwwx4 = (Yswwx4 & Ftwwx4);
assign Ftwwx4 = (~(hresp_i & H3owx4));
assign Yswwx4 = (Mtwwx4 & Ttwwx4);
assign Ttwwx4 = (~(Auwwx4 & G9lwx4));
assign G9lwx4 = (~(Huwwx4 & Ouwwx4));
assign Ouwwx4 = (~(hrdata_i[7] & B7owx4));
assign Huwwx4 = (Vuwwx4 & Cvwwx4);
assign Cvwwx4 = (~(L5owx4 & Fq7wx4));
assign Fq7wx4 = (Yw7wx4 ? Vzdwx4 : Nodwx4);
assign Vzdwx4 = (~(Jvwwx4 & Qvwwx4));
assign Qvwwx4 = (Xvwwx4 & Ewwwx4);
assign Ewwwx4 = (~(O1qwx4 & Niqwx4));
assign Xvwwx4 = (A1qwx4 | Ai9wx4);
assign Jvwwx4 = (Lwwwx4 & Swwwx4);
assign Swwwx4 = (~(Yzpwx4 & Wjqwx4));
assign Lwwwx4 = (~(Kzpwx4 & Uluwx4));
assign Nodwx4 = (~(Zwwwx4 & Gxwwx4));
assign Gxwwx4 = (Nxwwx4 & Uxwwx4);
assign Uxwwx4 = (~(O1qwx4 & Quqwx4));
assign Nxwwx4 = (A1qwx4 | Bywwx4);
assign Zwwwx4 = (Iywwx4 & Pywwx4);
assign Pywwx4 = (~(Yzpwx4 & Xuqwx4));
assign Iywwx4 = (~(Kzpwx4 & I0vwx4));
assign Vuwwx4 = (~(H3owx4 & Wywwx4));
assign Wywwx4 = (~(Dzwwx4 & Kzwwx4));
assign Kzwwx4 = (Rzwwx4 & Yzwwx4);
assign Yzwwx4 = (F0xwx4 & M0xwx4);
assign M0xwx4 = (E0uvx4 | T0xwx4);
assign F0xwx4 = (Qwowx4 | A1xwx4);
assign Rzwwx4 = (H1xwx4 & O1xwx4);
assign O1xwx4 = (K7pwx4 | V1xwx4);
assign H1xwx4 = (N1uvx4 | C2xwx4);
assign Dzwwx4 = (J2xwx4 & Q2xwx4);
assign Q2xwx4 = (X2xwx4 & E3xwx4);
assign E3xwx4 = (~(T1i2z4[7] & Ts5wx4));
assign X2xwx4 = (~(M5tvx4 & L0i2z4[7]));
assign J2xwx4 = (L3xwx4 & S3xwx4);
assign S3xwx4 = (~(Irh2z4[7] & Japwx4));
assign L3xwx4 = (~(Czh2z4[7] & H6tvx4));
assign Auwwx4 = (~(Y47wx4 & Z3xwx4));
assign Z3xwx4 = (~(G4xwx4 & W5yvx4));
assign G4xwx4 = (~(B1ovx4 & N4xwx4));
assign N4xwx4 = (Zph2z4[0] | Zph2z4[1]);
assign Y47wx4 = (!Zocwx4);
assign Mtwwx4 = (U4xwx4 | Sr2wx4);
assign U4xwx4 = (Ifnwx4 ? B5xwx4 : Dswwx4);
assign Ifnwx4 = (!Zph2z4[0]);
assign B5xwx4 = (~(Zph2z4[1] & Walwx4));
assign Walwx4 = (~(I5xwx4 & P5xwx4));
assign P5xwx4 = (W5xwx4 & D6xwx4);
assign D6xwx4 = (~(hrdata_i[23] & B7owx4));
assign W5xwx4 = (K6xwx4 & R6xwx4);
assign R6xwx4 = (~(H3owx4 & Y6xwx4));
assign Y6xwx4 = (~(F7xwx4 & M7xwx4));
assign M7xwx4 = (T7xwx4 & A8xwx4);
assign A8xwx4 = (Qwowx4 | H8xwx4);
assign T7xwx4 = (O8xwx4 & V8xwx4);
assign V8xwx4 = (K3uvx4 | C9xwx4);
assign O8xwx4 = (E0uvx4 | J9xwx4);
assign F7xwx4 = (Q9xwx4 & X9xwx4);
assign X9xwx4 = (K7pwx4 | Eaxwx4);
assign Q9xwx4 = (N1uvx4 | Laxwx4);
assign K6xwx4 = (Lcowx4 | Xs7wx4);
assign Xs7wx4 = (Oldwx4 ? Zaxwx4 : Saxwx4);
assign Zaxwx4 = (!Uvdwx4);
assign Uvdwx4 = (~(Gbxwx4 & Nbxwx4));
assign Nbxwx4 = (Ubxwx4 & Bcxwx4);
assign Bcxwx4 = (~(O1qwx4 & E3qwx4));
assign Ubxwx4 = (A1qwx4 | Icxwx4);
assign Gbxwx4 = (Pcxwx4 & Wcxwx4);
assign Wcxwx4 = (~(Yzpwx4 & L3qwx4));
assign Pcxwx4 = (~(Kzpwx4 & Z6uwx4));
assign Saxwx4 = (Yvtwx4 & Fwtwx4);
assign Fwtwx4 = (Ddxwx4 & Kdxwx4);
assign Kdxwx4 = (~(O1qwx4 & Ddqwx4));
assign Ddxwx4 = (~(Kzpwx4 & Zruwx4));
assign Yvtwx4 = (Rdxwx4 & Ydxwx4);
assign Ydxwx4 = (A1qwx4 | Fexwx4);
assign Rdxwx4 = (~(Yzpwx4 & Meqwx4));
assign I5xwx4 = (Mexwx4 & Texwx4);
assign Texwx4 = (~(Irh2z4[23] & I7owx4));
assign I7owx4 = (H3owx4 & Japwx4);
assign Mexwx4 = (~(G6owx4 & Czh2z4[23]));
assign G6owx4 = (H3owx4 & H6tvx4);
assign Dswwx4 = (!Afxwx4);
assign Afxwx4 = (N7nwx4 ? U9lwx4 : Palwx4);
assign N7nwx4 = (!Zph2z4[1]);
assign U9lwx4 = (~(Hfxwx4 & Ofxwx4));
assign Ofxwx4 = (~(hrdata_i[15] & B7owx4));
assign Hfxwx4 = (Vfxwx4 & Cgxwx4);
assign Cgxwx4 = (~(L5owx4 & Tq7wx4));
assign Tq7wx4 = (Oldwx4 ? X0ewx4 : Qtdwx4);
assign X0ewx4 = (~(Jgxwx4 & Qgxwx4));
assign Qgxwx4 = (Xgxwx4 & Ehxwx4);
assign Ehxwx4 = (~(O1qwx4 & Flqwx4));
assign Xgxwx4 = (A1qwx4 | Ey9wx4);
assign Jgxwx4 = (Lhxwx4 & Shxwx4);
assign Shxwx4 = (~(Yzpwx4 & Mlqwx4));
assign Lhxwx4 = (~(Kzpwx4 & Sduwx4));
assign Qtdwx4 = (~(Zhxwx4 & Gixwx4));
assign Gixwx4 = (Nixwx4 & Uixwx4);
assign Uixwx4 = (~(O1qwx4 & Rzpwx4));
assign Nixwx4 = (A1qwx4 | Bjxwx4);
assign Zhxwx4 = (Ijxwx4 & Pjxwx4);
assign Pjxwx4 = (~(Yzpwx4 & V1qwx4));
assign Ijxwx4 = (~(Kzpwx4 & Y9uwx4));
assign Vfxwx4 = (~(H3owx4 & Wjxwx4));
assign Wjxwx4 = (~(Dkxwx4 & Kkxwx4));
assign Kkxwx4 = (Rkxwx4 & Ykxwx4);
assign Ykxwx4 = (Flxwx4 & Mlxwx4);
assign Mlxwx4 = (Qwowx4 | Tlxwx4);
assign Flxwx4 = (Amxwx4 & X3pwx4);
assign X3pwx4 = (Hmxwx4 | Xahvx4);
assign Amxwx4 = (E0uvx4 | Omxwx4);
assign Rkxwx4 = (Vmxwx4 & Cnxwx4);
assign Cnxwx4 = (~(N4rvx4 & Gc4wx4));
assign Gc4wx4 = (!Wfuwx4);
assign N4rvx4 = (Q4owx4 & Jnxwx4);
assign Jnxwx4 = (~(Qnxwx4 & Qjuwx4));
assign Qjuwx4 = (!X4owx4);
assign Qnxwx4 = (~(I6pwx4 | E5owx4));
assign Q4owx4 = (!L4pwx4);
assign L4pwx4 = (~(Dguwx4 & Yguwx4));
assign Dguwx4 = (~(Krgvx4 | Eqgvx4));
assign Vmxwx4 = (K7pwx4 | Xnxwx4);
assign Dkxwx4 = (Eoxwx4 & Loxwx4);
assign Loxwx4 = (Soxwx4 & Zoxwx4);
assign Zoxwx4 = (~(M5tvx4 & L0i2z4[15]));
assign M5tvx4 = (Gpxwx4 & Npxwx4);
assign Soxwx4 = (Upxwx4 & Bqxwx4);
assign Bqxwx4 = (N1uvx4 | Iqxwx4);
assign Upxwx4 = (~(T1i2z4[15] & Ts5wx4));
assign Ts5wx4 = (Pqxwx4 & Npxwx4);
assign Eoxwx4 = (Wqxwx4 & Drxwx4);
assign Drxwx4 = (~(Irh2z4[15] & Japwx4));
assign Japwx4 = (!T4uvx4);
assign T4uvx4 = (~(Krxwx4 & G8twx4));
assign G8twx4 = (Rrxwx4 & B5hvx4);
assign Rrxwx4 = (~(N6hvx4 | Xahvx4));
assign Wqxwx4 = (~(Czh2z4[15] & H6tvx4));
assign H6tvx4 = (Yrxwx4 & Dotwx4);
assign Yrxwx4 = (Pqxwx4 & Aiovx4);
assign Palwx4 = (~(Fsxwx4 & Msxwx4));
assign Msxwx4 = (~(hrdata_i[31] & B7owx4));
assign B7owx4 = (Tsxwx4 & Vssvx4);
assign Vssvx4 = (Atxwx4 & Htxwx4);
assign Htxwx4 = (~(L9hvx4 | Xahvx4));
assign Atxwx4 = (~(B5hvx4 | N6hvx4));
assign Tsxwx4 = (~(Lstwx4 | Z7hvx4));
assign Fsxwx4 = (Otxwx4 & Vtxwx4);
assign Vtxwx4 = (~(L5owx4 & Hr7wx4));
assign Hr7wx4 = (Juxwx4 ? U2ewx4 : Cuxwx4);
assign Juxwx4 = (Quxwx4 & Wdpwx4);
assign Wdpwx4 = (~(M3ovx4 | C9qwx4));
assign C9qwx4 = (Xuxwx4 & Yw7wx4);
assign Quxwx4 = (Vpuwx4 ? Weowx4 : Udowx4);
assign Vpuwx4 = (!A1qwx4);
assign Weowx4 = (Yw7wx4 | Xuxwx4);
assign Udowx4 = (!Xuxwx4);
assign Xuxwx4 = (Dp7wx4 & Klwwx4);
assign Klwwx4 = (~(Evxwx4 & Dw7wx4));
assign Dw7wx4 = (Pkwwx4 & Vy7wx4);
assign Vy7wx4 = (F3ovx4 ? Svxwx4 : Lvxwx4);
assign Lvxwx4 = (~(Zvxwx4 & Vk7wx4));
assign Vk7wx4 = (~(Gwxwx4 & Svxwx4));
assign Zvxwx4 = (Svxwx4 | Gwxwx4);
assign Svxwx4 = (Nwxwx4 & Uwxwx4);
assign Uwxwx4 = (Bxxwx4 | Ixxwx4);
assign Nwxwx4 = (~(Hnwwx4 & Yo9vx4));
assign Pkwwx4 = (F3ovx4 ? Wxxwx4 : Pxxwx4);
assign Pxxwx4 = (Dyxwx4 | Gwxwx4);
assign Gwxwx4 = (Kyxwx4 & Wxxwx4);
assign Dyxwx4 = (~(Kyxwx4 | Wxxwx4));
assign Wxxwx4 = (Ryxwx4 & Yyxwx4);
assign Yyxwx4 = (Bxxwx4 | Fzxwx4);
assign Ryxwx4 = (~(Hnwwx4 & Un9vx4));
assign Kyxwx4 = (Mzxwx4 & Tzxwx4);
assign Evxwx4 = (~(Yw7wx4 | A1qwx4));
assign Yw7wx4 = (!Oldwx4);
assign Dp7wx4 = (!Z1ewx4);
assign Z1ewx4 = (~(Z6gvx4 | Eznvx4));
assign U2ewx4 = (A0ywx4 & Dw8vx4);
assign A0ywx4 = (H0ywx4 & Nbqwx4);
assign H0ywx4 = (~(O0ywx4 & Db7wx4));
assign O0ywx4 = (M93wx4 | Z6gvx4);
assign Cuxwx4 = (Oldwx4 ? Kw7wx4 : Rw7wx4);
assign Oldwx4 = (F3ovx4 ? Tzxwx4 : V0ywx4);
assign V0ywx4 = (~(Mzxwx4 ^ Tzxwx4));
assign Tzxwx4 = (C1ywx4 & J1ywx4);
assign J1ywx4 = (Bxxwx4 | Q1ywx4);
assign C1ywx4 = (~(Hnwwx4 & Qm9vx4));
assign Kw7wx4 = (~(X1ywx4 & E2ywx4));
assign E2ywx4 = (L2ywx4 & S2ywx4);
assign S2ywx4 = (~(O1qwx4 & Ubqwx4));
assign L2ywx4 = (~(Yzpwx4 & Laqwx4));
assign X1ywx4 = (Z2ywx4 & G3ywx4);
assign G3ywx4 = (A1qwx4 | N3ywx4);
assign Z2ywx4 = (~(Kzpwx4 & Ituwx4));
assign Rw7wx4 = (~(U3ywx4 & B4ywx4));
assign B4ywx4 = (I4ywx4 & P4ywx4);
assign P4ywx4 = (~(O1qwx4 & Bqqwx4));
assign O1qwx4 = (~(W4ywx4 | D5ywx4));
assign I4ywx4 = (~(Yzpwx4 & Drqwx4));
assign Yzpwx4 = (D5ywx4 & W4ywx4);
assign U3ywx4 = (K5ywx4 & R5ywx4);
assign R5ywx4 = (A1qwx4 | Ebbwx4);
assign A1qwx4 = (~(D5ywx4 & Y5ywx4));
assign K5ywx4 = (~(Kzpwx4 & Lyuwx4));
assign Kzpwx4 = (~(D5ywx4 | Y5ywx4));
assign D5ywx4 = (F3ovx4 ? M6ywx4 : F6ywx4);
assign F6ywx4 = (T6ywx4 | Mzxwx4);
assign Mzxwx4 = (~(A7ywx4 | W4ywx4));
assign T6ywx4 = (~(Y5ywx4 | M6ywx4));
assign M6ywx4 = (!A7ywx4);
assign A7ywx4 = (~(H7ywx4 & O7ywx4));
assign O7ywx4 = (Bxxwx4 | V7ywx4);
assign H7ywx4 = (~(Hnwwx4 & Ml9vx4));
assign Y5ywx4 = (!W4ywx4);
assign W4ywx4 = (~(C8ywx4 & J8ywx4));
assign J8ywx4 = (Bxxwx4 | Q8ywx4);
assign Bxxwx4 = (!Cowwx4);
assign Cowwx4 = (~(Ev5wx4 | F57wx4));
assign F57wx4 = (!Wkxvx4);
assign C8ywx4 = (~(Hnwwx4 & Ik9vx4));
assign Hnwwx4 = (Dw8vx4 & Sy2wx4);
assign L5owx4 = (!Lcowx4);
assign Lcowx4 = (~(Dw8vx4 & X8ywx4));
assign X8ywx4 = (~(E9ywx4 & L9ywx4));
assign L9ywx4 = (B1ovx4 | Ncqvx4);
assign E9ywx4 = (~(Locwx4 | Zocwx4));
assign Otxwx4 = (~(H3owx4 & S9ywx4));
assign S9ywx4 = (~(Z9ywx4 & Gaywx4));
assign Gaywx4 = (Naywx4 & Uaywx4);
assign Uaywx4 = (Bbywx4 & Ibywx4);
assign Ibywx4 = (~(P2uvx4 & Uth2z4[1]));
assign P2uvx4 = (Pbywx4 & Gpxwx4);
assign Bbywx4 = (K3uvx4 | Wbywx4);
assign K3uvx4 = (~(Krxwx4 & Dcywx4));
assign Dcywx4 = (Kcywx4 & N6hvx4);
assign Kcywx4 = (~(B5hvx4 | Xahvx4));
assign Krxwx4 = (~(Aiovx4 | Jjovx4));
assign Naywx4 = (Rcywx4 & Ycywx4);
assign Ycywx4 = (E0uvx4 | Fdywx4);
assign E0uvx4 = (Mdywx4 | Xahvx4);
assign Rcywx4 = (Qwowx4 | Tdywx4);
assign Qwowx4 = (Mdywx4 | Rgovx4);
assign Mdywx4 = (~(Aeywx4 & L9hvx4));
assign Aeywx4 = (Pqxwx4 & N6hvx4);
assign Pqxwx4 = (B5hvx4 & Jjovx4);
assign Z9ywx4 = (Heywx4 & Oeywx4);
assign Oeywx4 = (Veywx4 & Cfywx4);
assign Cfywx4 = (K7pwx4 | Jfywx4);
assign K7pwx4 = (Qfywx4 | Rgovx4);
assign Veywx4 = (N1uvx4 | Xfywx4);
assign N1uvx4 = (Qfywx4 | Xahvx4);
assign Qfywx4 = (~(Egywx4 & B5hvx4));
assign Egywx4 = (Z7hvx4 & Npxwx4);
assign Heywx4 = (Zipwx4 & Lgywx4);
assign Lgywx4 = (Sw4wx4 | Wfuwx4);
assign Wfuwx4 = (Rgovx4 | Hmxwx4);
assign Hmxwx4 = (~(Sgywx4 & Z7hvx4));
assign Sgywx4 = (Npxwx4 & X5ovx4);
assign Npxwx4 = (N6hvx4 & Aiovx4);
assign Zipwx4 = (~(Z4wwx4 | Zgywx4));
assign Zgywx4 = (Pbywx4 & Ghywx4);
assign Ghywx4 = (~(X5ovx4 | Jjovx4));
assign Jjovx4 = (!Z7hvx4);
assign X5ovx4 = (!B5hvx4);
assign Pbywx4 = (L9hvx4 & Dotwx4);
assign Dotwx4 = (Xahvx4 & Zkovx4);
assign Zkovx4 = (!N6hvx4);
assign Nqwwx4 = (~(Nhywx4 & Uhywx4));
assign Uhywx4 = (Biywx4 & W8nwx4);
assign W8nwx4 = (~(Iiywx4 & E6nwx4));
assign Iiywx4 = (hresp_i & H3owx4);
assign H3owx4 = (!Lstwx4);
assign Lstwx4 = (Ev5wx4 | Piywx4);
assign Piywx4 = (Wiywx4 & Djywx4);
assign Djywx4 = (B1ovx4 ? Kjywx4 : Agqvx4);
assign Kjywx4 = (Bdqvx4 | U0ovx4);
assign Agqvx4 = (!M5swx4);
assign M5swx4 = (~(S87wx4 | U9gvx4));
assign Wiywx4 = (Rjywx4 & Zrvvx4);
assign Rjywx4 = (Mvgwx4 | Cn8vx4);
assign Ev5wx4 = (!Dw8vx4);
assign Biywx4 = (~(Yjywx4 & Wdxvx4));
assign Yjywx4 = (~(Izwvx4 | Us2wx4));
assign Nhywx4 = (E6nwx4 & Fkywx4);
assign Fkywx4 = (~(Nggvx4 & Hw2wx4));
assign E6nwx4 = (~(Locwx4 | Mkywx4));
assign Mkywx4 = (Tkywx4 & Bdqvx4);
assign Tkywx4 = (~(Qaqvx4 | Fjgvx4));
assign Locwx4 = (~(Whgvx4 | Fjgvx4));
assign Lefwx4 = (~(G6pvx4 & Alywx4));
assign Alywx4 = (~(Hlywx4 & Olywx4));
assign Olywx4 = (~(Ul8vx4 & F3vvx4));
assign Hlywx4 = (Vlywx4 & Z5pvx4);
assign Vlywx4 = (~(Lrvvx4 & Mk8vx4));
assign Lrvvx4 = (~(Gxqvx4 | S6vvx4));
assign G6pvx4 = (!Qaiwx4);
assign Qaiwx4 = (~(hready_i & Dcrwx4));
assign Edhvx4 = (~(Cmywx4 & Jmywx4));
assign Jmywx4 = (~(H0gvx4 & Qmywx4));
assign Qmywx4 = (E7mwx4 | Ccovx4);
assign Cmywx4 = (Xmywx4 | Ccovx4);
assign Ccovx4 = (!hready_i);
assign Xchvx4 = (hready_i ? Enywx4 : Cvgvx4);
assign Enywx4 = (Lnywx4 & Snywx4);
assign Snywx4 = (Znywx4 & Goywx4);
assign Goywx4 = (~(Noywx4 & Ih8vx4));
assign Noywx4 = (Ffqvx4 & Ps3wx4);
assign Znywx4 = (~(Ki8vx4 & Uoywx4));
assign Uoywx4 = (~(Bpywx4 & Ipywx4));
assign Ipywx4 = (Sznvx4 | Us2wx4);
assign Bpywx4 = (Mu3wx4 | Vdgvx4);
assign Lnywx4 = (Abovx4 & Ppywx4);
assign Ppywx4 = (~(H8jwx4 & Pkiwx4));
assign Pkiwx4 = (M93wx4 | Ws3wx4);
assign Ws3wx4 = (Wpywx4 & Dqywx4);
assign Dqywx4 = (~(P5jwx4 & Clewx4));
assign P5jwx4 = (~(Mv2wx4 | Nggvx4));
assign Wpywx4 = (Yplwx4 | Whgvx4);
assign Yplwx4 = (~(Kqywx4 & Kngwx4));
assign Kqywx4 = (~(Mj8vx4 | Cn8vx4));
assign H8jwx4 = (Yt3wx4 | Us2wx4);
assign Abovx4 = (Rqywx4 & Yqywx4);
assign Yqywx4 = (~(Frywx4 & C6mwx4));
assign C6mwx4 = (Mrywx4 & Trywx4);
assign Trywx4 = (~(Asywx4 & Hsywx4));
assign Hsywx4 = (~(Osywx4 & Vsywx4));
assign Osywx4 = (E5owx4 ? Jtywx4 : Ctywx4);
assign Asywx4 = (Qtywx4 & Xtywx4);
assign Qtywx4 = (~(Euywx4 & Luywx4));
assign Euywx4 = (G5pwx4 ? Zuywx4 : Suywx4);
assign Zuywx4 = (Gvywx4 & Nvywx4);
assign Nvywx4 = (Vsywx4 | Ctywx4);
assign Suywx4 = (Uvywx4 & Bwywx4);
assign Bwywx4 = (Jtywx4 | Vsywx4);
assign Uvywx4 = (S4pwx4 ? Iwywx4 : Sxowx4);
assign Mrywx4 = (Yguwx4 & S6vvx4);
assign Yguwx4 = (~(Pwywx4 & G5pwx4));
assign G5pwx4 = (!E5owx4);
assign E5owx4 = (Wwywx4 & Dxywx4);
assign Dxywx4 = (~(Kxywx4 & Rxywx4));
assign Rxywx4 = (~(Yxywx4 & Fyywx4));
assign Fyywx4 = (~(Myywx4 & Tyywx4));
assign Tyywx4 = (S4pwx4 ? Uth2z4[0] : Psh2z4[0]);
assign Myywx4 = (Gvywx4 & Azywx4);
assign Azywx4 = (Ctywx4 | Hzywx4);
assign Ctywx4 = (!Ozywx4);
assign Gvywx4 = (C0zwx4 ? Vzywx4 : Vgpwx4);
assign Yxywx4 = (Jtywx4 | Ozywx4);
assign Ozywx4 = (C0zwx4 ? J0zwx4 : Txh2z4[1]);
assign Jtywx4 = (!Hzywx4);
assign Hzywx4 = (Avvwx4 ? Psh2z4[1] : Uth2z4[1]);
assign Avvwx4 = (!S4pwx4);
assign Kxywx4 = (~(X4owx4 & C0zwx4));
assign Wwywx4 = (Qsgvx4 | S4pwx4);
assign S4pwx4 = (Wtgvx4 & Q0zwx4);
assign Q0zwx4 = (~(X0zwx4 & Qsgvx4));
assign X0zwx4 = (E1zwx4 & L1zwx4);
assign L1zwx4 = (S1zwx4 | Uth2z4[1]);
assign S1zwx4 = (Z1zwx4 & C9xwx4);
assign E1zwx4 = (C9xwx4 | Z1zwx4);
assign Z1zwx4 = (~(Iwywx4 | Psh2z4[0]));
assign Pwywx4 = (X4owx4 & C0zwx4);
assign X4owx4 = (~(G2zwx4 & C0zwx4));
assign C0zwx4 = (~(R3hvx4 & N2zwx4));
assign N2zwx4 = (~(U2zwx4 & B3zwx4));
assign B3zwx4 = (~(J0zwx4 & Wbywx4));
assign U2zwx4 = (G2zwx4 & I3zwx4);
assign I3zwx4 = (~(P3zwx4 & W3zwx4));
assign W3zwx4 = (~(Vzywx4 & Txh2z4[0]));
assign Vzywx4 = (D4zwx4 & K4zwx4);
assign K4zwx4 = (I6pwx4 | R4zwx4);
assign D4zwx4 = (~(I6pwx4 & Y4zwx4));
assign Y4zwx4 = (~(F5zwx4 & M5zwx4));
assign F5zwx4 = (B6pwx4 | T5zwx4);
assign P3zwx4 = (J0zwx4 | Wbywx4);
assign J0zwx4 = (I6pwx4 ? H6zwx4 : A6zwx4);
assign G2zwx4 = (~(O6zwx4 & Hiuwx4));
assign O6zwx4 = (V6zwx4 & I6pwx4);
assign I6pwx4 = (~(C7zwx4 & J7zwx4));
assign J7zwx4 = (~(Q7zwx4 & X7zwx4));
assign X7zwx4 = (~(E8zwx4 & L8zwx4));
assign L8zwx4 = (~(S8zwx4 & Z8zwx4));
assign Z8zwx4 = (G9zwx4 & M5zwx4);
assign M5zwx4 = (~(B6pwx4 & N9zwx4));
assign N9zwx4 = (~(U9zwx4 & Bazwx4));
assign U9zwx4 = (Iazwx4 | Pazwx4);
assign G9zwx4 = (~(H6zwx4 & Wazwx4));
assign S8zwx4 = (~(R4zwx4 | Dbzwx4));
assign Dbzwx4 = (~(B6pwx4 | T5zwx4));
assign R4zwx4 = (U5pwx4 ? Rbzwx4 : Kbzwx4);
assign E8zwx4 = (Wazwx4 | H6zwx4);
assign H6zwx4 = (B6pwx4 ? Fczwx4 : Ybzwx4);
assign Ybzwx4 = (!Mczwx4);
assign Wazwx4 = (!A6zwx4);
assign A6zwx4 = (U5pwx4 ? Adzwx4 : Tczwx4);
assign Tczwx4 = (!Hdzwx4);
assign Q7zwx4 = (~(Hiuwx4 & V6zwx4));
assign Hiuwx4 = (B6pwx4 & Sxvwx4);
assign B6pwx4 = (~(Odzwx4 & Vdzwx4));
assign Vdzwx4 = (~(Cezwx4 & Jezwx4));
assign Cezwx4 = (~(Viuwx4 | Gyvwx4));
assign Odzwx4 = (~(Qezwx4 & Xezwx4));
assign Xezwx4 = (~(Efzwx4 & Lfzwx4));
assign Lfzwx4 = (~(Sfzwx4 & Zfzwx4));
assign Zfzwx4 = (Ggzwx4 & Bazwx4);
assign Bazwx4 = (~(Pazwx4 & Ngzwx4));
assign Ggzwx4 = (~(Fczwx4 & Mczwx4));
assign Sfzwx4 = (~(T5zwx4 | Ugzwx4));
assign Ugzwx4 = (~(Iazwx4 | Pazwx4));
assign T5zwx4 = (Phzwx4 ? Ihzwx4 : Bhzwx4);
assign Bhzwx4 = (Whzwx4 ? J3pwx4 : Tmpwx4);
assign Efzwx4 = (Mczwx4 | Fczwx4);
assign Fczwx4 = (Sxvwx4 ? Kizwx4 : Dizwx4);
assign Sxvwx4 = (!Pazwx4);
assign Mczwx4 = (Phzwx4 ? Yizwx4 : Rizwx4);
assign Phzwx4 = (!Viuwx4);
assign Viuwx4 = (Fjzwx4 & Mjzwx4);
assign Mjzwx4 = (~(Tjzwx4 & Akzwx4));
assign Akzwx4 = (~(Hkzwx4 & Okzwx4));
assign Okzwx4 = (~(Vkzwx4 & Clzwx4));
assign Clzwx4 = (Nyvwx4 ? Zuh2z4[16] : Zuh2z4[18]);
assign Nyvwx4 = (!Whzwx4);
assign Vkzwx4 = (Ihzwx4 & Jlzwx4);
assign Jlzwx4 = (Yizwx4 | Qlzwx4);
assign Ihzwx4 = (Gyvwx4 ? Zxowx4 : Chpwx4);
assign Hkzwx4 = (~(Qlzwx4 & Yizwx4));
assign Tjzwx4 = (~(Jezwx4 & Xlzwx4));
assign Fjzwx4 = (~(Whzwx4 & Emzwx4));
assign Emzwx4 = (~(T1i2z4[9] & L0i2z4[9]));
assign Yizwx4 = (Xlzwx4 ? Fdywx4 : J9xwx4);
assign Xlzwx4 = (!Gyvwx4);
assign Gyvwx4 = (Lmzwx4 & T1i2z4[10]);
assign Lmzwx4 = (L0i2z4[10] & Smzwx4);
assign Smzwx4 = (Jezwx4 | Zmzwx4);
assign Zmzwx4 = (Gnzwx4 & Nnzwx4);
assign Nnzwx4 = (~(Unzwx4 & Zuh2z4[20]));
assign Unzwx4 = (Bozwx4 & Chpwx4);
assign Bozwx4 = (Fdywx4 | Zuh2z4[21]);
assign Gnzwx4 = (J9xwx4 | Zuh2z4[23]);
assign Jezwx4 = (~(T1i2z4[11] & L0i2z4[11]));
assign Rizwx4 = (!Qlzwx4);
assign Qlzwx4 = (Whzwx4 ? Zuh2z4[19] : Zuh2z4[17]);
assign Whzwx4 = (~(Iozwx4 & T1i2z4[8]));
assign Iozwx4 = (L0i2z4[8] & Pozwx4);
assign Pozwx4 = (~(Wozwx4 & Dpzwx4));
assign Dpzwx4 = (Kpzwx4 & Rpzwx4);
assign Rpzwx4 = (~(Ypzwx4 & Fqzwx4));
assign Fqzwx4 = (T0xwx4 | Zuh2z4[19]);
assign Ypzwx4 = (Tmpwx4 | Zuh2z4[18]);
assign Kpzwx4 = (Omxwx4 | Zuh2z4[17]);
assign Wozwx4 = (T1i2z4[9] & L0i2z4[9]);
assign Qezwx4 = (Mqzwx4 | Pazwx4);
assign Pazwx4 = (Tqzwx4 & Arzwx4);
assign Arzwx4 = (~(Mqzwx4 & Hrzwx4));
assign Hrzwx4 = (~(Orzwx4 & Vrzwx4));
assign Vrzwx4 = (~(Cszwx4 & Ngzwx4));
assign Ngzwx4 = (Zxvwx4 ? Zuh2z4[24] : Zuh2z4[26]);
assign Cszwx4 = (Iazwx4 & Jszwx4);
assign Jszwx4 = (~(Qszwx4 & Kizwx4));
assign Iazwx4 = (Xwvwx4 ? Lipwx4 : Xwowx4);
assign Orzwx4 = (Kizwx4 | Qszwx4);
assign Qszwx4 = (!Dizwx4);
assign Dizwx4 = (Xszwx4 ? Zuh2z4[27] : Zuh2z4[25]);
assign Kizwx4 = (Xwvwx4 ? Zuh2z4[31] : Zuh2z4[29]);
assign Tqzwx4 = (~(Xszwx4 & Etzwx4));
assign Etzwx4 = (~(T1i2z4[13] & L0i2z4[13]));
assign Xszwx4 = (!Zxvwx4);
assign Zxvwx4 = (Ltzwx4 & T1i2z4[12]);
assign Ltzwx4 = (L0i2z4[12] & Stzwx4);
assign Stzwx4 = (~(Ztzwx4 & Guzwx4));
assign Guzwx4 = (Nuzwx4 & Uuzwx4);
assign Uuzwx4 = (~(Bvzwx4 & Ivzwx4));
assign Ivzwx4 = (A1xwx4 | Zuh2z4[27]);
assign Bvzwx4 = (~(Zuh2z4[24] & D7pwx4));
assign Nuzwx4 = (Tlxwx4 | Zuh2z4[25]);
assign Ztzwx4 = (T1i2z4[13] & L0i2z4[13]);
assign C7zwx4 = (~(Pvzwx4 & Wvzwx4));
assign Pvzwx4 = (Dwzwx4 & U5pwx4);
assign U5pwx4 = (~(Kwzwx4 & Rwzwx4));
assign Rwzwx4 = (~(Ywzwx4 & Fxzwx4));
assign Ywzwx4 = (~(Cjuwx4 | D0wwx4));
assign Kwzwx4 = (~(Mxzwx4 & Txzwx4));
assign Txzwx4 = (~(Wvzwx4 & Dwzwx4));
assign Wvzwx4 = (~(Jjuwx4 | Ayzwx4));
assign Mxzwx4 = (~(Hyzwx4 & Oyzwx4));
assign Oyzwx4 = (~(Vyzwx4 & Rbzwx4));
assign Rbzwx4 = (!Czzwx4);
assign Czzwx4 = (Xzzwx4 ? Qzzwx4 : Jzzwx4);
assign Vyzwx4 = (~(Kbzwx4 | E00xx4));
assign E00xx4 = (Adzwx4 & Hdzwx4);
assign Kbzwx4 = (Z00xx4 ? S00xx4 : L00xx4);
assign L00xx4 = (G10xx4 ? O9pwx4 : Onpwx4);
assign Hyzwx4 = (Hdzwx4 | Adzwx4);
assign Adzwx4 = (Xzzwx4 ? U10xx4 : N10xx4);
assign Xzzwx4 = (!Jjuwx4);
assign Jjuwx4 = (B20xx4 & I20xx4);
assign I20xx4 = (~(P20xx4 & W20xx4));
assign W20xx4 = (~(D30xx4 & K30xx4));
assign K30xx4 = (~(R30xx4 & Jzzwx4));
assign Jzzwx4 = (Wzvwx4 ? Zuh2z4[10] : Zuh2z4[8]);
assign R30xx4 = (~(Qzzwx4 | Y30xx4));
assign Y30xx4 = (~(F40xx4 | N10xx4));
assign Qzzwx4 = (Pzvwx4 ? Zuh2z4[14] : Zuh2z4[12]);
assign D30xx4 = (~(N10xx4 & F40xx4));
assign P20xx4 = (~(Dwzwx4 & Pzvwx4));
assign B20xx4 = (~(Wzvwx4 & M40xx4));
assign M40xx4 = (~(T1i2z4[5] & L0i2z4[5]));
assign U10xx4 = (!F40xx4);
assign F40xx4 = (Pzvwx4 ? Jfywx4 : Eaxwx4);
assign Pzvwx4 = (!Ayzwx4);
assign Ayzwx4 = (T40xx4 & T1i2z4[6]);
assign T40xx4 = (L0i2z4[6] & A50xx4);
assign A50xx4 = (H50xx4 | Dwzwx4);
assign H50xx4 = (~(O50xx4 & V50xx4));
assign V50xx4 = (~(C60xx4 & J60xx4));
assign J60xx4 = (Eaxwx4 | Zuh2z4[15]);
assign C60xx4 = (~(Zuh2z4[12] & Sipwx4));
assign O50xx4 = (Jfywx4 | Zuh2z4[13]);
assign N10xx4 = (Wzvwx4 ? Zuh2z4[11] : Zuh2z4[9]);
assign Wzvwx4 = (~(Q60xx4 & T1i2z4[4]));
assign Q60xx4 = (L0i2z4[4] & X60xx4);
assign X60xx4 = (~(E70xx4 & L70xx4));
assign L70xx4 = (S70xx4 & Z70xx4);
assign Z70xx4 = (~(G80xx4 & N80xx4));
assign N80xx4 = (V1xwx4 | Zuh2z4[11]);
assign G80xx4 = (~(Zuh2z4[8] & R7pwx4));
assign S70xx4 = (Xnxwx4 | Zuh2z4[9]);
assign E70xx4 = (T1i2z4[5] & L0i2z4[5]);
assign Hdzwx4 = (Z00xx4 ? B90xx4 : U80xx4);
assign Z00xx4 = (!Cjuwx4);
assign Cjuwx4 = (I90xx4 & P90xx4);
assign P90xx4 = (~(W90xx4 & Da0xx4));
assign Da0xx4 = (~(Ka0xx4 & Ra0xx4));
assign Ra0xx4 = (~(Ya0xx4 & Fb0xx4));
assign Fb0xx4 = (K0wwx4 ? Zuh2z4[0] : Zuh2z4[2]);
assign K0wwx4 = (!G10xx4);
assign Ya0xx4 = (S00xx4 & Mb0xx4);
assign Mb0xx4 = (B90xx4 | Tb0xx4);
assign S00xx4 = (D0wwx4 ? Uyowx4 : Njpwx4);
assign Ka0xx4 = (~(Tb0xx4 & B90xx4));
assign W90xx4 = (~(Fxzwx4 & Ac0xx4));
assign I90xx4 = (~(G10xx4 & Hc0xx4));
assign Hc0xx4 = (~(T1i2z4[1] & L0i2z4[1]));
assign B90xx4 = (Ac0xx4 ? Xfywx4 : Laxwx4);
assign Ac0xx4 = (!D0wwx4);
assign D0wwx4 = (Oc0xx4 & T1i2z4[2]);
assign Oc0xx4 = (L0i2z4[2] & Vc0xx4);
assign Vc0xx4 = (Fxzwx4 | Cd0xx4);
assign Cd0xx4 = (Jd0xx4 & Qd0xx4);
assign Qd0xx4 = (~(Xd0xx4 & Zuh2z4[4]));
assign Xd0xx4 = (Ee0xx4 & Njpwx4);
assign Ee0xx4 = (Xfywx4 | Zuh2z4[5]);
assign Jd0xx4 = (Laxwx4 | Zuh2z4[7]);
assign Fxzwx4 = (~(T1i2z4[3] & L0i2z4[3]));
assign U80xx4 = (!Tb0xx4);
assign Tb0xx4 = (G10xx4 ? Zuh2z4[3] : Zuh2z4[1]);
assign G10xx4 = (~(Le0xx4 & T1i2z4[0]));
assign Le0xx4 = (L0i2z4[0] & Se0xx4);
assign Se0xx4 = (~(Ze0xx4 & Gf0xx4));
assign Gf0xx4 = (Nf0xx4 & Uf0xx4);
assign Uf0xx4 = (~(Bg0xx4 & Ig0xx4));
assign Ig0xx4 = (C2xwx4 | Zuh2z4[3]);
assign Bg0xx4 = (Onpwx4 | Zuh2z4[2]);
assign Nf0xx4 = (Iqxwx4 | Zuh2z4[1]);
assign Ze0xx4 = (T1i2z4[1] & L0i2z4[1]);
assign Dwzwx4 = (~(T1i2z4[7] & L0i2z4[7]));
assign V6zwx4 = (!Mqzwx4);
assign Mqzwx4 = (~(Xwvwx4 & Pg0xx4));
assign Pg0xx4 = (~(T1i2z4[15] & L0i2z4[15]));
assign Xwvwx4 = (~(Wg0xx4 & T1i2z4[14]));
assign Wg0xx4 = (L0i2z4[14] & Dh0xx4);
assign Dh0xx4 = (~(Kh0xx4 & Rh0xx4));
assign Rh0xx4 = (Yh0xx4 & Fi0xx4);
assign Fi0xx4 = (~(Mi0xx4 & Ti0xx4));
assign Ti0xx4 = (H8xwx4 | Zuh2z4[31]);
assign Mi0xx4 = (Xwowx4 | Zuh2z4[30]);
assign Yh0xx4 = (Tdywx4 | Zuh2z4[29]);
assign Kh0xx4 = (T1i2z4[15] & L0i2z4[15]);
assign Frywx4 = (Gjqvx4 & Ujqvx4);
assign Ujqvx4 = (~(Aj0xx4 & Hj0xx4));
assign Hj0xx4 = (~(Oj0xx4 & Vj0xx4));
assign Vj0xx4 = (~(Ck0xx4 & B73wx4));
assign Ck0xx4 = (Z9dwx4 & Fs8vx4);
assign Oj0xx4 = (~(Kd5wx4 & Kryvx4));
assign Kd5wx4 = (!Zhyvx4);
assign Aj0xx4 = (Jk0xx4 | Qk0xx4);
assign Gjqvx4 = (~(Xk0xx4 & vis_primask_o));
assign Xk0xx4 = (~(Jk0xx4 | Qk0xx4));
assign Qk0xx4 = (El0xx4 & Yo9vx4);
assign El0xx4 = (Kryvx4 & Yryvx4);
assign Kryvx4 = (~(Ll0xx4 & Sl0xx4));
assign Sl0xx4 = (~(Zl0xx4 & Sy2wx4));
assign Zl0xx4 = (R13wx4 & W5yvx4);
assign Ll0xx4 = (Keqvx4 | M3ovx4);
assign Jk0xx4 = (Gm0xx4 & Nm0xx4);
assign Nm0xx4 = (~(S4xvx4 | Yg2wx4));
assign Yg2wx4 = (Um0xx4 & Bn0xx4);
assign Bn0xx4 = (Wm2wx4 & In0xx4);
assign In0xx4 = (~(Tjh2z4[1] & Qj2wx4));
assign Qj2wx4 = (~(Pn0xx4 & Wn0xx4));
assign Wn0xx4 = (Do0xx4 & Ko0xx4);
assign Ko0xx4 = (~(Ro0xx4 | Wbkwx4));
assign Wbkwx4 = (~(Fscwx4 | Efgvx4));
assign Ro0xx4 = (Yo0xx4 & Whgvx4);
assign Yo0xx4 = (Dbgvx4 & Fp0xx4);
assign Fp0xx4 = (~(Oedwx4 & Mp0xx4));
assign Mp0xx4 = (Vdgvx4 | Fjgvx4);
assign Do0xx4 = (Tp0xx4 & Aq0xx4);
assign Aq0xx4 = (~(Q43wx4 & Howvx4));
assign Q43wx4 = (~(U9gvx4 | Z6gvx4));
assign Tp0xx4 = (~(Wkxvx4 & Mcgvx4));
assign Pn0xx4 = (Hq0xx4 & Oq0xx4);
assign Oq0xx4 = (S4xvx4 ? Cr0xx4 : Vq0xx4);
assign Cr0xx4 = (M93wx4 | Nggvx4);
assign Vq0xx4 = (F3ovx4 | Bl3wx4);
assign Hq0xx4 = (Jucwx4 & Jr0xx4);
assign Jr0xx4 = (Gcqvx4 | Efgvx4);
assign Jucwx4 = (Hp2wx4 & Qr0xx4);
assign Qr0xx4 = (~(Wlhwx4 & Z7fwx4));
assign Wlhwx4 = (~(Gcqvx4 | O4ovx4));
assign Wm2wx4 = (~(Xr0xx4 | I7pvx4));
assign Xr0xx4 = (Es0xx4 & Nggvx4);
assign Es0xx4 = (Hw2wx4 & Izwvx4);
assign Um0xx4 = (Ls0xx4 & Ss0xx4);
assign Ss0xx4 = (~(Su9vx4 & Oi2wx4));
assign Oi2wx4 = (~(Zs0xx4 & Gt0xx4));
assign Gt0xx4 = (Zf7wx4 & Mu3wx4);
assign Mu3wx4 = (~(Nt0xx4 & O9qvx4));
assign Nt0xx4 = (~(M93wx4 | Nggvx4));
assign Zf7wx4 = (~(Wxcwx4 & Wkxvx4));
assign Zs0xx4 = (Ut0xx4 & Bu0xx4);
assign Bu0xx4 = (~(Iu0xx4 & Ncqvx4));
assign Iu0xx4 = (~(S4xvx4 | B1ovx4));
assign Ut0xx4 = (~(Cn8vx4 & Pu0xx4));
assign Pu0xx4 = (~(Wu0xx4 & Lbqvx4));
assign Lbqvx4 = (Zj3wx4 | U9gvx4);
assign Wu0xx4 = (Dv0xx4 & Kv0xx4);
assign Kv0xx4 = (~(Z9dwx4 & Nggvx4));
assign Dv0xx4 = (Tv2wx4 | U0ovx4);
assign Ls0xx4 = (~(Fs8vx4 & Vi2wx4));
assign Vi2wx4 = (~(Rv0xx4 & Yv0xx4));
assign Yv0xx4 = (Njxvx4 | Us2wx4);
assign Rv0xx4 = (Fw0xx4 & Mw0xx4);
assign Mw0xx4 = (~(Tw0xx4 & Z3jwx4));
assign Z3jwx4 = (~(U0ovx4 | Bl3wx4));
assign Tw0xx4 = (~(B4dwx4 | Bdqvx4));
assign Bdqvx4 = (!Y13wx4);
assign B4dwx4 = (!Ax0xx4);
assign Fw0xx4 = (~(Hx0xx4 & Ox0xx4));
assign Ox0xx4 = (~(Cn8vx4 | Z6gvx4));
assign Hx0xx4 = (~(Gcqvx4 | Mvgwx4));
assign Gm0xx4 = (B73wx4 & Z9dwx4);
assign Rqywx4 = (Q6mwx4 | F3vvx4);
assign F3vvx4 = (~(S6vvx4 | vis_ipsr_o[0]));
assign S6vvx4 = (!Ye4wx4);
assign Q6mwx4 = (Sw4wx4 & Vx0xx4);
assign Vx0xx4 = (Ytvwx4 | Ye4wx4);
assign Ytvwx4 = (!Krgvx4);
assign Sw4wx4 = (!Eqgvx4);
assign Qchvx4 = (~(Jchvx4 & Cy0xx4));
assign Cy0xx4 = (~(Jy0xx4 & Qy0xx4));
assign Qy0xx4 = (Xy0xx4 & Ez0xx4);
assign Ez0xx4 = (Lz0xx4 & Sz0xx4);
assign Sz0xx4 = (D04wx4 & Sx3wx4);
assign D04wx4 = (~(hwdata_o[29] | hwdata_o[30]));
assign hwdata_o[30] = (~(Zz0xx4 & G01xx4));
assign G01xx4 = (~(N01xx4 & El8wx4));
assign El8wx4 = (!S71wx4);
assign S71wx4 = (U01xx4 & B11xx4);
assign B11xx4 = (I11xx4 & P11xx4);
assign P11xx4 = (W11xx4 & D21xx4);
assign D21xx4 = (K21xx4 & R21xx4);
assign R21xx4 = (~(vis_psp_o[12] & Y21xx4));
assign K21xx4 = (F31xx4 & M31xx4);
assign M31xx4 = (~(vis_r6_o[14] & T31xx4));
assign F31xx4 = (~(vis_r0_o[14] & A41xx4));
assign W11xx4 = (H41xx4 & O41xx4);
assign O41xx4 = (~(vis_r1_o[14] & V41xx4));
assign H41xx4 = (~(vis_msp_o[12] & C51xx4));
assign I11xx4 = (J51xx4 & Q51xx4);
assign Q51xx4 = (X51xx4 & E61xx4);
assign E61xx4 = (~(vis_r14_o[14] & L61xx4));
assign X51xx4 = (~(vis_r2_o[14] & S61xx4));
assign J51xx4 = (Z61xx4 & G71xx4);
assign G71xx4 = (~(vis_r12_o[14] & N71xx4));
assign Z61xx4 = (~(vis_r5_o[14] & U71xx4));
assign U01xx4 = (B81xx4 & I81xx4);
assign I81xx4 = (P81xx4 & W81xx4);
assign W81xx4 = (D91xx4 & K91xx4);
assign K91xx4 = (~(vis_r4_o[14] & R91xx4));
assign D91xx4 = (~(vis_r11_o[14] & Y91xx4));
assign P81xx4 = (Fa1xx4 & Ma1xx4);
assign Ma1xx4 = (~(Yhdvx4 & Ta1xx4));
assign Fa1xx4 = (~(vis_r9_o[14] & Ab1xx4));
assign B81xx4 = (Hb1xx4 & Ob1xx4);
assign Ob1xx4 = (Vb1xx4 & Cc1xx4);
assign Cc1xx4 = (~(vis_r7_o[14] & Jc1xx4));
assign Vb1xx4 = (~(vis_r3_o[14] & Qc1xx4));
assign Hb1xx4 = (Xc1xx4 & Ed1xx4);
assign Ed1xx4 = (~(vis_r10_o[14] & Ld1xx4));
assign Xc1xx4 = (~(vis_r8_o[14] & Sd1xx4));
assign Zz0xx4 = (Zd1xx4 & Pq5wx4);
assign Pq5wx4 = (Yd5wx4 | Uvzvx4);
assign Zd1xx4 = (~(Ge1xx4 & H2bwx4));
assign H2bwx4 = (!O7zvx4);
assign O7zvx4 = (Ne1xx4 & Ue1xx4);
assign Ue1xx4 = (Bf1xx4 & If1xx4);
assign If1xx4 = (Pf1xx4 & Wf1xx4);
assign Wf1xx4 = (Dg1xx4 & Kg1xx4);
assign Kg1xx4 = (~(S4evx4 & Ta1xx4));
assign Dg1xx4 = (Rg1xx4 & Yg1xx4);
assign Yg1xx4 = (~(vis_psp_o[28] & Y21xx4));
assign Rg1xx4 = (~(vis_msp_o[28] & C51xx4));
assign Pf1xx4 = (Fh1xx4 & Mh1xx4);
assign Mh1xx4 = (~(vis_r14_o[30] & L61xx4));
assign Fh1xx4 = (~(vis_r12_o[30] & N71xx4));
assign Bf1xx4 = (Th1xx4 & Ai1xx4);
assign Ai1xx4 = (Hi1xx4 & Oi1xx4);
assign Oi1xx4 = (~(vis_r11_o[30] & Y91xx4));
assign Hi1xx4 = (~(vis_r10_o[30] & Ld1xx4));
assign Th1xx4 = (Vi1xx4 & Cj1xx4);
assign Cj1xx4 = (~(vis_r9_o[30] & Ab1xx4));
assign Vi1xx4 = (~(vis_r8_o[30] & Sd1xx4));
assign Ne1xx4 = (Jj1xx4 & Qj1xx4);
assign Qj1xx4 = (Xj1xx4 & Ek1xx4);
assign Ek1xx4 = (Lk1xx4 & Sk1xx4);
assign Sk1xx4 = (~(vis_r7_o[30] & Jc1xx4));
assign Lk1xx4 = (~(vis_r6_o[30] & T31xx4));
assign Xj1xx4 = (Zk1xx4 & Gl1xx4);
assign Gl1xx4 = (~(vis_r5_o[30] & U71xx4));
assign Zk1xx4 = (~(vis_r4_o[30] & R91xx4));
assign Jj1xx4 = (Nl1xx4 & Ul1xx4);
assign Ul1xx4 = (Bm1xx4 & Im1xx4);
assign Im1xx4 = (~(vis_r3_o[30] & Qc1xx4));
assign Bm1xx4 = (~(vis_r2_o[30] & S61xx4));
assign Nl1xx4 = (Pm1xx4 & Wm1xx4);
assign Wm1xx4 = (~(vis_r1_o[30] & V41xx4));
assign Pm1xx4 = (~(vis_r0_o[30] & A41xx4));
assign Lz0xx4 = (~(hwdata_o[25] | hwdata_o[27]));
assign Xy0xx4 = (Dn1xx4 & Kn1xx4);
assign Kn1xx4 = (hwdata_o[26] & Ux4wx4);
assign Ux4wx4 = (~(Mf8vx4 & hwdata_o[31]));
assign Dn1xx4 = (~(hwdata_o[18] | Rn1xx4));
assign Rn1xx4 = (!hwdata_o[24]);
assign hwdata_o[18] = (Ge1xx4 ? Aj8wx4 : Sh5wx4);
assign Aj8wx4 = (!St0wx4);
assign St0wx4 = (Yn1xx4 & Fo1xx4);
assign Fo1xx4 = (Mo1xx4 & To1xx4);
assign To1xx4 = (Ap1xx4 & Hp1xx4);
assign Hp1xx4 = (Op1xx4 & Vp1xx4);
assign Vp1xx4 = (~(Qndvx4 & Ta1xx4));
assign Op1xx4 = (Cq1xx4 & Jq1xx4);
assign Jq1xx4 = (~(vis_psp_o[16] & Y21xx4));
assign Cq1xx4 = (~(vis_msp_o[16] & C51xx4));
assign Ap1xx4 = (Qq1xx4 & Xq1xx4);
assign Xq1xx4 = (~(vis_r14_o[18] & L61xx4));
assign Qq1xx4 = (~(vis_r12_o[18] & N71xx4));
assign Mo1xx4 = (Er1xx4 & Lr1xx4);
assign Lr1xx4 = (Sr1xx4 & Zr1xx4);
assign Zr1xx4 = (~(vis_r11_o[18] & Y91xx4));
assign Sr1xx4 = (~(vis_r10_o[18] & Ld1xx4));
assign Er1xx4 = (Gs1xx4 & Ns1xx4);
assign Ns1xx4 = (~(vis_r9_o[18] & Ab1xx4));
assign Gs1xx4 = (~(vis_r8_o[18] & Sd1xx4));
assign Yn1xx4 = (Us1xx4 & Bt1xx4);
assign Bt1xx4 = (It1xx4 & Pt1xx4);
assign Pt1xx4 = (Wt1xx4 & Du1xx4);
assign Du1xx4 = (~(vis_r7_o[18] & Jc1xx4));
assign Wt1xx4 = (~(vis_r6_o[18] & T31xx4));
assign It1xx4 = (Ku1xx4 & Ru1xx4);
assign Ru1xx4 = (~(vis_r5_o[18] & U71xx4));
assign Ku1xx4 = (~(vis_r4_o[18] & R91xx4));
assign Us1xx4 = (Yu1xx4 & Fv1xx4);
assign Fv1xx4 = (Mv1xx4 & Tv1xx4);
assign Tv1xx4 = (~(vis_r3_o[18] & Qc1xx4));
assign Mv1xx4 = (~(vis_r2_o[18] & S61xx4));
assign Yu1xx4 = (Aw1xx4 & Hw1xx4);
assign Hw1xx4 = (~(vis_r1_o[18] & V41xx4));
assign Aw1xx4 = (~(vis_r0_o[18] & A41xx4));
assign Jy0xx4 = (Ow1xx4 & Vw1xx4);
assign Vw1xx4 = (Cx1xx4 & Jx1xx4);
assign Jx1xx4 = (Qx1xx4 & Z4wwx4);
assign Z4wwx4 = (Xx1xx4 & Ey1xx4);
assign Ey1xx4 = (Gpxwx4 & N6hvx4);
assign Gpxwx4 = (~(B5hvx4 | Z7hvx4));
assign Xx1xx4 = (~(Aiovx4 | Rgovx4));
assign Rgovx4 = (!Xahvx4);
assign Aiovx4 = (!L9hvx4);
assign Qx1xx4 = (V4ovx4 & O24wx4);
assign O24wx4 = (Ge1xx4 ? W21wx4 : Zhyvx4);
assign W21wx4 = (Ly1xx4 & Sy1xx4);
assign Sy1xx4 = (Zy1xx4 & Gz1xx4);
assign Gz1xx4 = (Nz1xx4 & Uz1xx4);
assign Uz1xx4 = (B02xx4 & I02xx4);
assign I02xx4 = (~(Ukdvx4 & Ta1xx4));
assign B02xx4 = (P02xx4 & W02xx4);
assign W02xx4 = (~(vis_psp_o[14] & Y21xx4));
assign P02xx4 = (~(vis_msp_o[14] & C51xx4));
assign Nz1xx4 = (D12xx4 & K12xx4);
assign K12xx4 = (~(vis_r14_o[16] & L61xx4));
assign D12xx4 = (~(vis_r12_o[16] & N71xx4));
assign Zy1xx4 = (R12xx4 & Y12xx4);
assign Y12xx4 = (F22xx4 & M22xx4);
assign M22xx4 = (~(vis_r11_o[16] & Y91xx4));
assign F22xx4 = (~(vis_r10_o[16] & Ld1xx4));
assign R12xx4 = (T22xx4 & A32xx4);
assign A32xx4 = (~(vis_r9_o[16] & Ab1xx4));
assign T22xx4 = (~(vis_r8_o[16] & Sd1xx4));
assign Ly1xx4 = (H32xx4 & O32xx4);
assign O32xx4 = (V32xx4 & C42xx4);
assign C42xx4 = (J42xx4 & Q42xx4);
assign Q42xx4 = (~(vis_r7_o[16] & Jc1xx4));
assign J42xx4 = (~(vis_r6_o[16] & T31xx4));
assign V32xx4 = (X42xx4 & E52xx4);
assign E52xx4 = (~(vis_r5_o[16] & U71xx4));
assign X42xx4 = (~(vis_r4_o[16] & R91xx4));
assign H32xx4 = (L52xx4 & S52xx4);
assign S52xx4 = (Z52xx4 & G62xx4);
assign G62xx4 = (~(vis_r3_o[16] & Qc1xx4));
assign Z52xx4 = (~(vis_r2_o[16] & S61xx4));
assign L52xx4 = (N62xx4 & U62xx4);
assign U62xx4 = (~(vis_r1_o[16] & V41xx4));
assign N62xx4 = (~(vis_r0_o[16] & A41xx4));
assign V4ovx4 = (Mf8vx4 & hwdata_o[23]);
assign Cx1xx4 = (hwdata_o[17] & hwdata_o[2]);
assign hwdata_o[2] = (!L35wx4);
assign L35wx4 = (~(Pp8vx4 & Sh5wx4));
assign hwdata_o[17] = (Ge1xx4 ? Hj8wx4 : Htyvx4);
assign Hj8wx4 = (!Yw0wx4);
assign Yw0wx4 = (B72xx4 & I72xx4);
assign I72xx4 = (P72xx4 & W72xx4);
assign W72xx4 = (D82xx4 & K82xx4);
assign K82xx4 = (R82xx4 & Y82xx4);
assign Y82xx4 = (~(Fmdvx4 & Ta1xx4));
assign R82xx4 = (F92xx4 & M92xx4);
assign M92xx4 = (~(vis_psp_o[15] & Y21xx4));
assign F92xx4 = (~(vis_msp_o[15] & C51xx4));
assign D82xx4 = (T92xx4 & Aa2xx4);
assign Aa2xx4 = (~(vis_r14_o[17] & L61xx4));
assign T92xx4 = (~(vis_r12_o[17] & N71xx4));
assign P72xx4 = (Ha2xx4 & Oa2xx4);
assign Oa2xx4 = (Va2xx4 & Cb2xx4);
assign Cb2xx4 = (~(vis_r11_o[17] & Y91xx4));
assign Va2xx4 = (~(vis_r10_o[17] & Ld1xx4));
assign Ha2xx4 = (Jb2xx4 & Qb2xx4);
assign Qb2xx4 = (~(vis_r9_o[17] & Ab1xx4));
assign Jb2xx4 = (~(vis_r8_o[17] & Sd1xx4));
assign B72xx4 = (Xb2xx4 & Ec2xx4);
assign Ec2xx4 = (Lc2xx4 & Sc2xx4);
assign Sc2xx4 = (Zc2xx4 & Gd2xx4);
assign Gd2xx4 = (~(vis_r7_o[17] & Jc1xx4));
assign Zc2xx4 = (~(vis_r6_o[17] & T31xx4));
assign Lc2xx4 = (Nd2xx4 & Ud2xx4);
assign Ud2xx4 = (~(vis_r5_o[17] & U71xx4));
assign Nd2xx4 = (~(vis_r4_o[17] & R91xx4));
assign Xb2xx4 = (Be2xx4 & Ie2xx4);
assign Ie2xx4 = (Pe2xx4 & We2xx4);
assign We2xx4 = (~(vis_r3_o[17] & Qc1xx4));
assign Pe2xx4 = (~(vis_r2_o[17] & S61xx4));
assign Be2xx4 = (Df2xx4 & Kf2xx4);
assign Kf2xx4 = (~(vis_r1_o[17] & V41xx4));
assign Df2xx4 = (~(vis_r0_o[17] & A41xx4));
assign Ow1xx4 = (Rf2xx4 & Yf2xx4);
assign Yf2xx4 = (hwdata_o[19] & hwdata_o[20]);
assign hwdata_o[20] = (Ge1xx4 ? Fg2xx4 : Am5wx4);
assign Fg2xx4 = (!Hk0wx4);
assign Hk0wx4 = (Mg2xx4 & Tg2xx4);
assign Tg2xx4 = (Ah2xx4 & Hh2xx4);
assign Hh2xx4 = (Oh2xx4 & Vh2xx4);
assign Vh2xx4 = (Ci2xx4 & Ji2xx4);
assign Ji2xx4 = (~(Mqdvx4 & Ta1xx4));
assign Ci2xx4 = (Qi2xx4 & Xi2xx4);
assign Xi2xx4 = (~(vis_psp_o[18] & Y21xx4));
assign Qi2xx4 = (~(vis_msp_o[18] & C51xx4));
assign Oh2xx4 = (Ej2xx4 & Lj2xx4);
assign Lj2xx4 = (~(vis_r14_o[20] & L61xx4));
assign Ej2xx4 = (~(vis_r12_o[20] & N71xx4));
assign Ah2xx4 = (Sj2xx4 & Zj2xx4);
assign Zj2xx4 = (Gk2xx4 & Nk2xx4);
assign Nk2xx4 = (~(vis_r11_o[20] & Y91xx4));
assign Gk2xx4 = (~(vis_r10_o[20] & Ld1xx4));
assign Sj2xx4 = (Uk2xx4 & Bl2xx4);
assign Bl2xx4 = (~(vis_r9_o[20] & Ab1xx4));
assign Uk2xx4 = (~(vis_r8_o[20] & Sd1xx4));
assign Mg2xx4 = (Il2xx4 & Pl2xx4);
assign Pl2xx4 = (Wl2xx4 & Dm2xx4);
assign Dm2xx4 = (Km2xx4 & Rm2xx4);
assign Rm2xx4 = (~(vis_r7_o[20] & Jc1xx4));
assign Km2xx4 = (~(vis_r6_o[20] & T31xx4));
assign Wl2xx4 = (Ym2xx4 & Fn2xx4);
assign Fn2xx4 = (~(vis_r5_o[20] & U71xx4));
assign Ym2xx4 = (~(vis_r4_o[20] & R91xx4));
assign Il2xx4 = (Mn2xx4 & Tn2xx4);
assign Tn2xx4 = (Ao2xx4 & Ho2xx4);
assign Ho2xx4 = (~(vis_r3_o[20] & Qc1xx4));
assign Ao2xx4 = (~(vis_r2_o[20] & S61xx4));
assign Mn2xx4 = (Oo2xx4 & Vo2xx4);
assign Vo2xx4 = (~(vis_r1_o[20] & V41xx4));
assign Oo2xx4 = (~(vis_r0_o[20] & A41xx4));
assign hwdata_o[19] = (Ge1xx4 ? Xk8wx4 : Wj5wx4);
assign Xk8wx4 = (!Nn0wx4);
assign Nn0wx4 = (Cp2xx4 & Jp2xx4);
assign Jp2xx4 = (Qp2xx4 & Xp2xx4);
assign Xp2xx4 = (Eq2xx4 & Lq2xx4);
assign Lq2xx4 = (Sq2xx4 & Zq2xx4);
assign Zq2xx4 = (~(Bpdvx4 & Ta1xx4));
assign Sq2xx4 = (Gr2xx4 & Nr2xx4);
assign Nr2xx4 = (~(vis_psp_o[17] & Y21xx4));
assign Gr2xx4 = (~(vis_msp_o[17] & C51xx4));
assign Eq2xx4 = (Ur2xx4 & Bs2xx4);
assign Bs2xx4 = (~(vis_r14_o[19] & L61xx4));
assign Ur2xx4 = (~(vis_r12_o[19] & N71xx4));
assign Qp2xx4 = (Is2xx4 & Ps2xx4);
assign Ps2xx4 = (Ws2xx4 & Dt2xx4);
assign Dt2xx4 = (~(vis_r11_o[19] & Y91xx4));
assign Ws2xx4 = (~(vis_r10_o[19] & Ld1xx4));
assign Is2xx4 = (Kt2xx4 & Rt2xx4);
assign Rt2xx4 = (~(vis_r9_o[19] & Ab1xx4));
assign Kt2xx4 = (~(vis_r8_o[19] & Sd1xx4));
assign Cp2xx4 = (Yt2xx4 & Fu2xx4);
assign Fu2xx4 = (Mu2xx4 & Tu2xx4);
assign Tu2xx4 = (Av2xx4 & Hv2xx4);
assign Hv2xx4 = (~(vis_r7_o[19] & Jc1xx4));
assign Av2xx4 = (~(vis_r6_o[19] & T31xx4));
assign Mu2xx4 = (Ov2xx4 & Vv2xx4);
assign Vv2xx4 = (~(vis_r5_o[19] & U71xx4));
assign Ov2xx4 = (~(vis_r4_o[19] & R91xx4));
assign Yt2xx4 = (Cw2xx4 & Jw2xx4);
assign Jw2xx4 = (Qw2xx4 & Xw2xx4);
assign Xw2xx4 = (~(vis_r3_o[19] & Qc1xx4));
assign Qw2xx4 = (~(vis_r2_o[19] & S61xx4));
assign Cw2xx4 = (Ex2xx4 & Lx2xx4);
assign Lx2xx4 = (~(vis_r1_o[19] & V41xx4));
assign Ex2xx4 = (~(vis_r0_o[19] & A41xx4));
assign Wj5wx4 = (!R40wx4);
assign Rf2xx4 = (hwdata_o[22] & hwdata_o[21]);
assign hwdata_o[21] = (Ge1xx4 ? Vj8wx4 : Eo5wx4);
assign Vj8wx4 = (!Ce0wx4);
assign Ce0wx4 = (Sx2xx4 & Zx2xx4);
assign Zx2xx4 = (Gy2xx4 & Ny2xx4);
assign Ny2xx4 = (Uy2xx4 & Bz2xx4);
assign Bz2xx4 = (Iz2xx4 & Pz2xx4);
assign Pz2xx4 = (~(Xrdvx4 & Ta1xx4));
assign Iz2xx4 = (Wz2xx4 & D03xx4);
assign D03xx4 = (~(vis_psp_o[19] & Y21xx4));
assign Wz2xx4 = (~(vis_msp_o[19] & C51xx4));
assign Uy2xx4 = (K03xx4 & R03xx4);
assign R03xx4 = (~(vis_r14_o[21] & L61xx4));
assign K03xx4 = (~(vis_r12_o[21] & N71xx4));
assign Gy2xx4 = (Y03xx4 & F13xx4);
assign F13xx4 = (M13xx4 & T13xx4);
assign T13xx4 = (~(vis_r11_o[21] & Y91xx4));
assign M13xx4 = (~(vis_r10_o[21] & Ld1xx4));
assign Y03xx4 = (A23xx4 & H23xx4);
assign H23xx4 = (~(vis_r9_o[21] & Ab1xx4));
assign A23xx4 = (~(vis_r8_o[21] & Sd1xx4));
assign Sx2xx4 = (O23xx4 & V23xx4);
assign V23xx4 = (C33xx4 & J33xx4);
assign J33xx4 = (Q33xx4 & X33xx4);
assign X33xx4 = (~(vis_r7_o[21] & Jc1xx4));
assign Q33xx4 = (~(vis_r6_o[21] & T31xx4));
assign C33xx4 = (E43xx4 & L43xx4);
assign L43xx4 = (~(vis_r5_o[21] & U71xx4));
assign E43xx4 = (~(vis_r4_o[21] & R91xx4));
assign O23xx4 = (S43xx4 & Z43xx4);
assign Z43xx4 = (G53xx4 & N53xx4);
assign N53xx4 = (~(vis_r3_o[21] & Qc1xx4));
assign G53xx4 = (~(vis_r2_o[21] & S61xx4));
assign S43xx4 = (U53xx4 & B63xx4);
assign B63xx4 = (~(vis_r1_o[21] & V41xx4));
assign U53xx4 = (~(vis_r0_o[21] & A41xx4));
assign hwdata_o[22] = (Ge1xx4 ? Qk8wx4 : Ll8wx4);
assign Qk8wx4 = (!Wa0wx4);
assign Wa0wx4 = (I63xx4 & P63xx4);
assign P63xx4 = (W63xx4 & D73xx4);
assign D73xx4 = (K73xx4 & R73xx4);
assign R73xx4 = (Y73xx4 & F83xx4);
assign F83xx4 = (~(Itdvx4 & Ta1xx4));
assign Y73xx4 = (M83xx4 & T83xx4);
assign T83xx4 = (~(vis_psp_o[20] & Y21xx4));
assign M83xx4 = (~(vis_msp_o[20] & C51xx4));
assign K73xx4 = (A93xx4 & H93xx4);
assign H93xx4 = (~(vis_r14_o[22] & L61xx4));
assign A93xx4 = (~(vis_r12_o[22] & N71xx4));
assign W63xx4 = (O93xx4 & V93xx4);
assign V93xx4 = (Ca3xx4 & Ja3xx4);
assign Ja3xx4 = (~(vis_r11_o[22] & Y91xx4));
assign Ca3xx4 = (~(vis_r10_o[22] & Ld1xx4));
assign O93xx4 = (Qa3xx4 & Xa3xx4);
assign Xa3xx4 = (~(vis_r9_o[22] & Ab1xx4));
assign Qa3xx4 = (~(vis_r8_o[22] & Sd1xx4));
assign I63xx4 = (Eb3xx4 & Lb3xx4);
assign Lb3xx4 = (Sb3xx4 & Zb3xx4);
assign Zb3xx4 = (Gc3xx4 & Nc3xx4);
assign Nc3xx4 = (~(vis_r7_o[22] & Jc1xx4));
assign Gc3xx4 = (~(vis_r6_o[22] & T31xx4));
assign Sb3xx4 = (Uc3xx4 & Bd3xx4);
assign Bd3xx4 = (~(vis_r5_o[22] & U71xx4));
assign Uc3xx4 = (~(vis_r4_o[22] & R91xx4));
assign Eb3xx4 = (Id3xx4 & Pd3xx4);
assign Pd3xx4 = (Wd3xx4 & De3xx4);
assign De3xx4 = (~(vis_r3_o[22] & Qc1xx4));
assign Wd3xx4 = (~(vis_r2_o[22] & S61xx4));
assign Id3xx4 = (Ke3xx4 & Re3xx4);
assign Re3xx4 = (~(vis_r1_o[22] & V41xx4));
assign Ke3xx4 = (~(vis_r0_o[22] & A41xx4));
assign Ll8wx4 = (!Uvzvx4);
assign lockup_o = (!Z5pvx4);
assign hwdata_o[7] = (!Youvx4);
assign Youvx4 = (~(Pp8vx4 & Ht5wx4));
assign hwdata_o[6] = (~(C5vvx4 | Uvzvx4));
assign Uvzvx4 = (Ye3xx4 & Ff3xx4);
assign Ff3xx4 = (Mf3xx4 & Tf3xx4);
assign Tf3xx4 = (Ag3xx4 & Hg3xx4);
assign Hg3xx4 = (~(vis_r11_o[6] & Y91xx4));
assign Ag3xx4 = (Og3xx4 & Vg3xx4);
assign Vg3xx4 = (~(vis_r9_o[6] & Ab1xx4));
assign Og3xx4 = (~(S6dvx4 & Ta1xx4));
assign Mf3xx4 = (Ch3xx4 & Jh3xx4);
assign Jh3xx4 = (~(vis_r10_o[6] & Ld1xx4));
assign Ch3xx4 = (~(vis_psp_o[4] & Y21xx4));
assign Ye3xx4 = (Qh3xx4 & Xh3xx4);
assign Xh3xx4 = (Ei3xx4 & Li3xx4);
assign Li3xx4 = (~(vis_r12_o[6] & N71xx4));
assign Ei3xx4 = (Si3xx4 & Zi3xx4);
assign Zi3xx4 = (~(vis_msp_o[4] & C51xx4));
assign Si3xx4 = (~(vis_r14_o[6] & L61xx4));
assign Qh3xx4 = (Qowwx4 & Gj3xx4);
assign Gj3xx4 = (~(vis_r8_o[6] & Sd1xx4));
assign Qowwx4 = (Nj3xx4 & Uj3xx4);
assign Uj3xx4 = (Bk3xx4 & Ik3xx4);
assign Ik3xx4 = (Pk3xx4 & Wk3xx4);
assign Wk3xx4 = (~(vis_r0_o[6] & A41xx4));
assign Pk3xx4 = (~(vis_r2_o[6] & S61xx4));
assign Bk3xx4 = (Dl3xx4 & Kl3xx4);
assign Kl3xx4 = (~(vis_r5_o[6] & U71xx4));
assign Dl3xx4 = (~(vis_r4_o[6] & R91xx4));
assign Nj3xx4 = (Rl3xx4 & Yl3xx4);
assign Yl3xx4 = (Fm3xx4 & Mm3xx4);
assign Mm3xx4 = (~(vis_r7_o[6] & Jc1xx4));
assign Fm3xx4 = (~(vis_r3_o[6] & Qc1xx4));
assign Rl3xx4 = (Tm3xx4 & An3xx4);
assign An3xx4 = (~(vis_r1_o[6] & V41xx4));
assign Tm3xx4 = (~(vis_r6_o[6] & T31xx4));
assign hwdata_o[5] = (!Dvuvx4);
assign Dvuvx4 = (~(Pp8vx4 & Eo5wx4));
assign hwdata_o[4] = (!Jyuvx4);
assign Jyuvx4 = (~(Pp8vx4 & Am5wx4));
assign hwdata_o[3] = (~(C5vvx4 | R40wx4));
assign hwdata_o[31] = (~(Hn3xx4 & On3xx4));
assign On3xx4 = (~(Wq5wx4 & Ht5wx4));
assign Hn3xx4 = (Vn3xx4 & Co3xx4);
assign Co3xx4 = (~(Ge1xx4 & Grawx4));
assign Grawx4 = (!Nd3wx4);
assign Nd3wx4 = (Jo3xx4 & Qo3xx4);
assign Qo3xx4 = (Xo3xx4 & Ep3xx4);
assign Ep3xx4 = (Lp3xx4 & Sp3xx4);
assign Sp3xx4 = (Zp3xx4 & Gq3xx4);
assign Gq3xx4 = (~(D6evx4 & Ta1xx4));
assign Zp3xx4 = (Nq3xx4 & Uq3xx4);
assign Uq3xx4 = (~(vis_psp_o[29] & Y21xx4));
assign Nq3xx4 = (~(vis_msp_o[29] & C51xx4));
assign Lp3xx4 = (Br3xx4 & Ir3xx4);
assign Ir3xx4 = (~(vis_r14_o[31] & L61xx4));
assign Br3xx4 = (~(vis_r12_o[31] & N71xx4));
assign Xo3xx4 = (Pr3xx4 & Wr3xx4);
assign Wr3xx4 = (Ds3xx4 & Ks3xx4);
assign Ks3xx4 = (~(vis_r11_o[31] & Y91xx4));
assign Ds3xx4 = (~(vis_r10_o[31] & Ld1xx4));
assign Pr3xx4 = (Rs3xx4 & Ys3xx4);
assign Ys3xx4 = (~(vis_r9_o[31] & Ab1xx4));
assign Rs3xx4 = (~(vis_r8_o[31] & Sd1xx4));
assign Jo3xx4 = (Ft3xx4 & Mt3xx4);
assign Mt3xx4 = (Tt3xx4 & Au3xx4);
assign Au3xx4 = (Hu3xx4 & Ou3xx4);
assign Ou3xx4 = (~(vis_r7_o[31] & Jc1xx4));
assign Hu3xx4 = (~(vis_r6_o[31] & T31xx4));
assign Tt3xx4 = (Vu3xx4 & Cv3xx4);
assign Cv3xx4 = (~(vis_r5_o[31] & U71xx4));
assign Vu3xx4 = (~(vis_r4_o[31] & R91xx4));
assign Ft3xx4 = (Jv3xx4 & Qv3xx4);
assign Qv3xx4 = (Xv3xx4 & Ew3xx4);
assign Ew3xx4 = (~(vis_r3_o[31] & Qc1xx4));
assign Xv3xx4 = (~(vis_r2_o[31] & S61xx4));
assign Jv3xx4 = (Lw3xx4 & Sw3xx4);
assign Sw3xx4 = (~(vis_r1_o[31] & V41xx4));
assign Lw3xx4 = (~(vis_r0_o[31] & A41xx4));
assign Vn3xx4 = (~(N01xx4 & Ot5wx4));
assign Ot5wx4 = (!Z62wx4);
assign Z62wx4 = (Zw3xx4 & Gx3xx4);
assign Gx3xx4 = (Nx3xx4 & Ux3xx4);
assign Ux3xx4 = (By3xx4 & Iy3xx4);
assign Iy3xx4 = (Py3xx4 & Wy3xx4);
assign Wy3xx4 = (~(vis_r6_o[15] & T31xx4));
assign Py3xx4 = (Dz3xx4 & Kz3xx4);
assign Kz3xx4 = (~(Jjdvx4 & Ta1xx4));
assign Dz3xx4 = (~(vis_r2_o[15] & S61xx4));
assign By3xx4 = (Rz3xx4 & Yz3xx4);
assign Yz3xx4 = (~(vis_r5_o[15] & U71xx4));
assign Rz3xx4 = (~(vis_r4_o[15] & R91xx4));
assign Nx3xx4 = (F04xx4 & M04xx4);
assign M04xx4 = (T04xx4 & A14xx4);
assign A14xx4 = (~(vis_r10_o[15] & Ld1xx4));
assign T04xx4 = (~(vis_psp_o[13] & Y21xx4));
assign F04xx4 = (H14xx4 & O14xx4);
assign O14xx4 = (~(vis_msp_o[13] & C51xx4));
assign H14xx4 = (~(vis_r14_o[15] & L61xx4));
assign Zw3xx4 = (V14xx4 & C24xx4);
assign C24xx4 = (J24xx4 & Q24xx4);
assign Q24xx4 = (X24xx4 & E34xx4);
assign E34xx4 = (~(vis_r12_o[15] & N71xx4));
assign X24xx4 = (~(vis_r9_o[15] & Ab1xx4));
assign J24xx4 = (L34xx4 & S34xx4);
assign S34xx4 = (~(vis_r8_o[15] & Sd1xx4));
assign L34xx4 = (~(vis_r1_o[15] & V41xx4));
assign V14xx4 = (Z34xx4 & G44xx4);
assign G44xx4 = (N44xx4 & U44xx4);
assign U44xx4 = (~(vis_r0_o[15] & A41xx4));
assign N44xx4 = (~(vis_r3_o[15] & Qc1xx4));
assign Z34xx4 = (B54xx4 & I54xx4);
assign I54xx4 = (~(vis_r7_o[15] & Jc1xx4));
assign B54xx4 = (~(vis_r11_o[15] & Y91xx4));
assign hwdata_o[29] = (~(P54xx4 & W54xx4));
assign W54xx4 = (~(N01xx4 & Lo5wx4));
assign Lo5wx4 = (!Hc1wx4);
assign Hc1wx4 = (D64xx4 & K64xx4);
assign K64xx4 = (R64xx4 & Y64xx4);
assign Y64xx4 = (F74xx4 & M74xx4);
assign M74xx4 = (T74xx4 & A84xx4);
assign A84xx4 = (~(vis_r6_o[13] & T31xx4));
assign T74xx4 = (H84xx4 & O84xx4);
assign O84xx4 = (~(Ngdvx4 & Ta1xx4));
assign H84xx4 = (~(vis_r2_o[13] & S61xx4));
assign F74xx4 = (V84xx4 & C94xx4);
assign C94xx4 = (~(vis_r5_o[13] & U71xx4));
assign V84xx4 = (~(vis_r4_o[13] & R91xx4));
assign R64xx4 = (J94xx4 & Q94xx4);
assign Q94xx4 = (X94xx4 & Ea4xx4);
assign Ea4xx4 = (~(vis_r10_o[13] & Ld1xx4));
assign X94xx4 = (~(vis_psp_o[11] & Y21xx4));
assign J94xx4 = (La4xx4 & Sa4xx4);
assign Sa4xx4 = (~(vis_msp_o[11] & C51xx4));
assign La4xx4 = (~(vis_r14_o[13] & L61xx4));
assign D64xx4 = (Za4xx4 & Gb4xx4);
assign Gb4xx4 = (Nb4xx4 & Ub4xx4);
assign Ub4xx4 = (Bc4xx4 & Ic4xx4);
assign Ic4xx4 = (~(vis_r12_o[13] & N71xx4));
assign Bc4xx4 = (~(vis_r9_o[13] & Ab1xx4));
assign Nb4xx4 = (Pc4xx4 & Wc4xx4);
assign Wc4xx4 = (~(vis_r8_o[13] & Sd1xx4));
assign Pc4xx4 = (~(vis_r1_o[13] & V41xx4));
assign Za4xx4 = (Dd4xx4 & Kd4xx4);
assign Kd4xx4 = (Rd4xx4 & Yd4xx4);
assign Yd4xx4 = (~(vis_r0_o[13] & A41xx4));
assign Rd4xx4 = (~(vis_r3_o[13] & Qc1xx4));
assign Dd4xx4 = (Fe4xx4 & Me4xx4);
assign Me4xx4 = (~(vis_r7_o[13] & Jc1xx4));
assign Fe4xx4 = (~(vis_r11_o[13] & Y91xx4));
assign P54xx4 = (Te4xx4 & Af4xx4);
assign Af4xx4 = (~(Wq5wx4 & Eo5wx4));
assign Eo5wx4 = (~(Hf4xx4 & Of4xx4));
assign Of4xx4 = (Vf4xx4 & Cg4xx4);
assign Cg4xx4 = (Jg4xx4 & Spwwx4);
assign Spwwx4 = (Qg4xx4 & Xg4xx4);
assign Xg4xx4 = (~(vis_r3_o[5] & Qc1xx4));
assign Qg4xx4 = (~(vis_r7_o[5] & Jc1xx4));
assign Jg4xx4 = (Eh4xx4 & Lh4xx4);
assign Lh4xx4 = (~(vis_psp_o[3] & Y21xx4));
assign Eh4xx4 = (~(vis_msp_o[3] & C51xx4));
assign Vf4xx4 = (Sh4xx4 & Zh4xx4);
assign Zh4xx4 = (~(vis_r12_o[5] & N71xx4));
assign Sh4xx4 = (Gi4xx4 & Ni4xx4);
assign Ni4xx4 = (~(I5dvx4 & Ta1xx4));
assign Gi4xx4 = (~(vis_r14_o[5] & L61xx4));
assign Hf4xx4 = (Ui4xx4 & Bj4xx4);
assign Bj4xx4 = (Ij4xx4 & Pj4xx4);
assign Pj4xx4 = (~(vis_r9_o[5] & Ab1xx4));
assign Ij4xx4 = (Wj4xx4 & Dk4xx4);
assign Dk4xx4 = (~(vis_r11_o[5] & Y91xx4));
assign Wj4xx4 = (~(vis_r10_o[5] & Ld1xx4));
assign Ui4xx4 = (Kk4xx4 & Zpwwx4);
assign Zpwwx4 = (Rk4xx4 & Yk4xx4);
assign Yk4xx4 = (~(vis_r0_o[5] & A41xx4));
assign Rk4xx4 = (~(vis_r1_o[5] & V41xx4));
assign Kk4xx4 = (Gqwwx4 & Fl4xx4);
assign Fl4xx4 = (~(vis_r8_o[5] & Sd1xx4));
assign Gqwwx4 = (Ml4xx4 & Tl4xx4);
assign Tl4xx4 = (Am4xx4 & Hm4xx4);
assign Hm4xx4 = (~(vis_r2_o[5] & S61xx4));
assign Am4xx4 = (~(vis_r5_o[5] & U71xx4));
assign Ml4xx4 = (Om4xx4 & Vm4xx4);
assign Vm4xx4 = (~(vis_r4_o[5] & R91xx4));
assign Om4xx4 = (~(vis_r6_o[5] & T31xx4));
assign Te4xx4 = (~(Ge1xx4 & Shcwx4));
assign Shcwx4 = (!Rtpvx4);
assign Rtpvx4 = (Cn4xx4 & Jn4xx4);
assign Jn4xx4 = (Qn4xx4 & Xn4xx4);
assign Xn4xx4 = (Eo4xx4 & Lo4xx4);
assign Lo4xx4 = (So4xx4 & Zo4xx4);
assign Zo4xx4 = (~(H3evx4 & Ta1xx4));
assign So4xx4 = (Gp4xx4 & Np4xx4);
assign Np4xx4 = (~(vis_psp_o[27] & Y21xx4));
assign Gp4xx4 = (~(vis_msp_o[27] & C51xx4));
assign Eo4xx4 = (Up4xx4 & Bq4xx4);
assign Bq4xx4 = (~(vis_r14_o[29] & L61xx4));
assign Up4xx4 = (~(vis_r12_o[29] & N71xx4));
assign Qn4xx4 = (Iq4xx4 & Pq4xx4);
assign Pq4xx4 = (Wq4xx4 & Dr4xx4);
assign Dr4xx4 = (~(vis_r11_o[29] & Y91xx4));
assign Wq4xx4 = (~(vis_r10_o[29] & Ld1xx4));
assign Iq4xx4 = (Kr4xx4 & Rr4xx4);
assign Rr4xx4 = (~(vis_r9_o[29] & Ab1xx4));
assign Kr4xx4 = (~(vis_r8_o[29] & Sd1xx4));
assign Cn4xx4 = (Yr4xx4 & Fs4xx4);
assign Fs4xx4 = (Ms4xx4 & Ts4xx4);
assign Ts4xx4 = (At4xx4 & Ht4xx4);
assign Ht4xx4 = (~(vis_r7_o[29] & Jc1xx4));
assign At4xx4 = (~(vis_r6_o[29] & T31xx4));
assign Ms4xx4 = (Ot4xx4 & Vt4xx4);
assign Vt4xx4 = (~(vis_r5_o[29] & U71xx4));
assign Ot4xx4 = (~(vis_r4_o[29] & R91xx4));
assign Yr4xx4 = (Cu4xx4 & Ju4xx4);
assign Ju4xx4 = (Qu4xx4 & Xu4xx4);
assign Xu4xx4 = (~(vis_r3_o[29] & Qc1xx4));
assign Qu4xx4 = (~(vis_r2_o[29] & S61xx4));
assign Cu4xx4 = (Ev4xx4 & Lv4xx4);
assign Lv4xx4 = (~(vis_r1_o[29] & V41xx4));
assign Ev4xx4 = (~(vis_r0_o[29] & A41xx4));
assign hwdata_o[28] = (!Sx3wx4);
assign Sx3wx4 = (Sv4xx4 & Zv4xx4);
assign Zv4xx4 = (~(N01xx4 & Hm5wx4));
assign Hm5wx4 = (!Ze1wx4);
assign Ze1wx4 = (Gw4xx4 & Nw4xx4);
assign Nw4xx4 = (Uw4xx4 & Bx4xx4);
assign Bx4xx4 = (Ix4xx4 & Px4xx4);
assign Px4xx4 = (Wx4xx4 & Dy4xx4);
assign Dy4xx4 = (~(vis_psp_o[10] & Y21xx4));
assign Wx4xx4 = (Ky4xx4 & Ry4xx4);
assign Ry4xx4 = (~(vis_r6_o[12] & T31xx4));
assign Ky4xx4 = (~(vis_r0_o[12] & A41xx4));
assign Ix4xx4 = (Yy4xx4 & Fz4xx4);
assign Fz4xx4 = (~(vis_r1_o[12] & V41xx4));
assign Yy4xx4 = (~(vis_msp_o[10] & C51xx4));
assign Uw4xx4 = (Mz4xx4 & Tz4xx4);
assign Tz4xx4 = (A05xx4 & H05xx4);
assign H05xx4 = (~(vis_r14_o[12] & L61xx4));
assign A05xx4 = (~(vis_r2_o[12] & S61xx4));
assign Mz4xx4 = (O05xx4 & V05xx4);
assign V05xx4 = (~(vis_r12_o[12] & N71xx4));
assign O05xx4 = (~(vis_r5_o[12] & U71xx4));
assign Gw4xx4 = (C15xx4 & J15xx4);
assign J15xx4 = (Q15xx4 & X15xx4);
assign X15xx4 = (E25xx4 & L25xx4);
assign L25xx4 = (~(vis_r4_o[12] & R91xx4));
assign E25xx4 = (~(vis_r11_o[12] & Y91xx4));
assign Q15xx4 = (S25xx4 & Z25xx4);
assign Z25xx4 = (~(Cfdvx4 & Ta1xx4));
assign S25xx4 = (~(vis_r9_o[12] & Ab1xx4));
assign C15xx4 = (G35xx4 & N35xx4);
assign N35xx4 = (U35xx4 & B45xx4);
assign B45xx4 = (~(vis_r7_o[12] & Jc1xx4));
assign U35xx4 = (~(vis_r3_o[12] & Qc1xx4));
assign G35xx4 = (I45xx4 & P45xx4);
assign P45xx4 = (~(vis_r10_o[12] & Ld1xx4));
assign I45xx4 = (~(vis_r8_o[12] & Sd1xx4));
assign Sv4xx4 = (W45xx4 & D55xx4);
assign D55xx4 = (~(Wq5wx4 & Am5wx4));
assign Am5wx4 = (~(K55xx4 & R55xx4));
assign R55xx4 = (Y55xx4 & F65xx4);
assign F65xx4 = (M65xx4 & T65xx4);
assign T65xx4 = (~(Y3dvx4 & Ta1xx4));
assign M65xx4 = (A75xx4 & H75xx4);
assign H75xx4 = (~(vis_psp_o[2] & Y21xx4));
assign A75xx4 = (~(vis_msp_o[2] & C51xx4));
assign Y55xx4 = (O75xx4 & V75xx4);
assign V75xx4 = (~(vis_r14_o[4] & L61xx4));
assign O75xx4 = (~(vis_r12_o[4] & N71xx4));
assign K55xx4 = (C85xx4 & J85xx4);
assign J85xx4 = (Q85xx4 & X85xx4);
assign X85xx4 = (~(vis_r9_o[4] & Ab1xx4));
assign Q85xx4 = (E95xx4 & L95xx4);
assign L95xx4 = (~(vis_r11_o[4] & Y91xx4));
assign E95xx4 = (~(vis_r10_o[4] & Ld1xx4));
assign C85xx4 = (Ixxwx4 & S95xx4);
assign S95xx4 = (~(vis_r8_o[4] & Sd1xx4));
assign Ixxwx4 = (Z95xx4 & Ga5xx4);
assign Ga5xx4 = (Na5xx4 & Ua5xx4);
assign Ua5xx4 = (Bb5xx4 & Ib5xx4);
assign Ib5xx4 = (~(vis_r7_o[4] & Jc1xx4));
assign Bb5xx4 = (~(vis_r6_o[4] & T31xx4));
assign Na5xx4 = (Pb5xx4 & Wb5xx4);
assign Wb5xx4 = (~(vis_r5_o[4] & U71xx4));
assign Pb5xx4 = (~(vis_r4_o[4] & R91xx4));
assign Z95xx4 = (Dc5xx4 & Kc5xx4);
assign Kc5xx4 = (Rc5xx4 & Yc5xx4);
assign Yc5xx4 = (~(vis_r3_o[4] & Qc1xx4));
assign Rc5xx4 = (~(vis_r2_o[4] & S61xx4));
assign Dc5xx4 = (Fd5xx4 & Md5xx4);
assign Md5xx4 = (~(vis_r1_o[4] & V41xx4));
assign Fd5xx4 = (~(vis_r0_o[4] & A41xx4));
assign W45xx4 = (~(Ge1xx4 & Aoawx4));
assign Aoawx4 = (!Izpvx4);
assign Izpvx4 = (Td5xx4 & Ae5xx4);
assign Ae5xx4 = (He5xx4 & Oe5xx4);
assign Oe5xx4 = (Ve5xx4 & Cf5xx4);
assign Cf5xx4 = (Jf5xx4 & Qf5xx4);
assign Qf5xx4 = (~(W1evx4 & Ta1xx4));
assign Jf5xx4 = (Xf5xx4 & Eg5xx4);
assign Eg5xx4 = (~(vis_psp_o[26] & Y21xx4));
assign Xf5xx4 = (~(vis_msp_o[26] & C51xx4));
assign Ve5xx4 = (Lg5xx4 & Sg5xx4);
assign Sg5xx4 = (~(vis_r14_o[28] & L61xx4));
assign Lg5xx4 = (~(vis_r12_o[28] & N71xx4));
assign He5xx4 = (Zg5xx4 & Gh5xx4);
assign Gh5xx4 = (Nh5xx4 & Uh5xx4);
assign Uh5xx4 = (~(vis_r11_o[28] & Y91xx4));
assign Nh5xx4 = (~(vis_r10_o[28] & Ld1xx4));
assign Zg5xx4 = (Bi5xx4 & Ii5xx4);
assign Ii5xx4 = (~(vis_r9_o[28] & Ab1xx4));
assign Bi5xx4 = (~(vis_r8_o[28] & Sd1xx4));
assign Td5xx4 = (Pi5xx4 & Wi5xx4);
assign Wi5xx4 = (Dj5xx4 & Kj5xx4);
assign Kj5xx4 = (Rj5xx4 & Yj5xx4);
assign Yj5xx4 = (~(vis_r7_o[28] & Jc1xx4));
assign Rj5xx4 = (~(vis_r6_o[28] & T31xx4));
assign Dj5xx4 = (Fk5xx4 & Mk5xx4);
assign Mk5xx4 = (~(vis_r5_o[28] & U71xx4));
assign Fk5xx4 = (~(vis_r4_o[28] & R91xx4));
assign Pi5xx4 = (Tk5xx4 & Al5xx4);
assign Al5xx4 = (Hl5xx4 & Ol5xx4);
assign Ol5xx4 = (~(vis_r3_o[28] & Qc1xx4));
assign Hl5xx4 = (~(vis_r2_o[28] & S61xx4));
assign Tk5xx4 = (Vl5xx4 & Cm5xx4);
assign Cm5xx4 = (~(vis_r1_o[28] & V41xx4));
assign Vl5xx4 = (~(vis_r0_o[28] & A41xx4));
assign hwdata_o[27] = (~(Jm5xx4 & Qm5xx4));
assign Qm5xx4 = (~(N01xx4 & Dk5wx4));
assign Dk5wx4 = (!Gm1wx4);
assign Gm1wx4 = (Xm5xx4 & En5xx4);
assign En5xx4 = (Ln5xx4 & Sn5xx4);
assign Sn5xx4 = (Zn5xx4 & Go5xx4);
assign Go5xx4 = (No5xx4 & Uo5xx4);
assign Uo5xx4 = (~(vis_psp_o[9] & Y21xx4));
assign No5xx4 = (Bp5xx4 & Ip5xx4);
assign Ip5xx4 = (~(vis_r6_o[11] & T31xx4));
assign Bp5xx4 = (~(vis_r0_o[11] & A41xx4));
assign Zn5xx4 = (Pp5xx4 & Wp5xx4);
assign Wp5xx4 = (~(vis_r1_o[11] & V41xx4));
assign Pp5xx4 = (~(vis_msp_o[9] & C51xx4));
assign Ln5xx4 = (Dq5xx4 & Kq5xx4);
assign Kq5xx4 = (Rq5xx4 & Yq5xx4);
assign Yq5xx4 = (~(vis_r14_o[11] & L61xx4));
assign Rq5xx4 = (~(vis_r2_o[11] & S61xx4));
assign Dq5xx4 = (Fr5xx4 & Mr5xx4);
assign Mr5xx4 = (~(vis_r12_o[11] & N71xx4));
assign Fr5xx4 = (~(vis_r5_o[11] & U71xx4));
assign Xm5xx4 = (Tr5xx4 & As5xx4);
assign As5xx4 = (Hs5xx4 & Os5xx4);
assign Os5xx4 = (Vs5xx4 & Ct5xx4);
assign Ct5xx4 = (~(vis_r4_o[11] & R91xx4));
assign Vs5xx4 = (~(vis_r11_o[11] & Y91xx4));
assign Hs5xx4 = (Jt5xx4 & Qt5xx4);
assign Qt5xx4 = (~(Rddvx4 & Ta1xx4));
assign Jt5xx4 = (~(vis_r9_o[11] & Ab1xx4));
assign Tr5xx4 = (Xt5xx4 & Eu5xx4);
assign Eu5xx4 = (Lu5xx4 & Su5xx4);
assign Su5xx4 = (~(vis_r7_o[11] & Jc1xx4));
assign Lu5xx4 = (~(vis_r3_o[11] & Qc1xx4));
assign Xt5xx4 = (Zu5xx4 & Gv5xx4);
assign Gv5xx4 = (~(vis_r10_o[11] & Ld1xx4));
assign Zu5xx4 = (~(vis_r8_o[11] & Sd1xx4));
assign Jm5xx4 = (Nv5xx4 & Uv5xx4);
assign Uv5xx4 = (Yd5wx4 | R40wx4);
assign R40wx4 = (Bw5xx4 & Iw5xx4);
assign Iw5xx4 = (Pw5xx4 & Ww5xx4);
assign Ww5xx4 = (Dx5xx4 & Ol22z4);
assign Ol22z4 = (~(vis_r11_o[3] & Y91xx4));
assign Dx5xx4 = (Vl22z4 & Cm22z4);
assign Cm22z4 = (~(vis_r9_o[3] & Ab1xx4));
assign Vl22z4 = (~(O2dvx4 & Ta1xx4));
assign Pw5xx4 = (Jm22z4 & Qm22z4);
assign Qm22z4 = (~(vis_r10_o[3] & Ld1xx4));
assign Jm22z4 = (~(vis_psp_o[1] & Y21xx4));
assign Bw5xx4 = (Xm22z4 & En22z4);
assign En22z4 = (Ln22z4 & Sn22z4);
assign Sn22z4 = (~(vis_r12_o[3] & N71xx4));
assign Ln22z4 = (Zn22z4 & Go22z4);
assign Go22z4 = (~(vis_msp_o[1] & C51xx4));
assign Zn22z4 = (~(vis_r14_o[3] & L61xx4));
assign Xm22z4 = (Fzxwx4 & No22z4);
assign No22z4 = (~(vis_r8_o[3] & Sd1xx4));
assign Fzxwx4 = (Uo22z4 & Bp22z4);
assign Bp22z4 = (Ip22z4 & Pp22z4);
assign Pp22z4 = (Wp22z4 & Dq22z4);
assign Dq22z4 = (~(vis_r2_o[3] & S61xx4));
assign Wp22z4 = (~(vis_r6_o[3] & T31xx4));
assign Ip22z4 = (Kq22z4 & Rq22z4);
assign Rq22z4 = (~(vis_r5_o[3] & U71xx4));
assign Kq22z4 = (~(vis_r4_o[3] & R91xx4));
assign Uo22z4 = (Yq22z4 & Fr22z4);
assign Fr22z4 = (Mr22z4 & Tr22z4);
assign Tr22z4 = (~(vis_r1_o[3] & V41xx4));
assign Mr22z4 = (~(vis_r0_o[3] & A41xx4));
assign Yq22z4 = (As22z4 & Hs22z4);
assign Hs22z4 = (~(vis_r3_o[3] & Qc1xx4));
assign As22z4 = (~(vis_r7_o[3] & Jc1xx4));
assign Nv5xx4 = (~(Ge1xx4 & Ucbwx4));
assign Ucbwx4 = (!Pdbwx4);
assign Pdbwx4 = (Os22z4 & Vs22z4);
assign Vs22z4 = (Ct22z4 & Jt22z4);
assign Jt22z4 = (Qt22z4 & Xt22z4);
assign Xt22z4 = (Eu22z4 & Lu22z4);
assign Lu22z4 = (~(L0evx4 & Ta1xx4));
assign Eu22z4 = (Su22z4 & Zu22z4);
assign Zu22z4 = (~(vis_psp_o[25] & Y21xx4));
assign Su22z4 = (~(vis_msp_o[25] & C51xx4));
assign Qt22z4 = (Gv22z4 & Nv22z4);
assign Nv22z4 = (~(vis_r14_o[27] & L61xx4));
assign Gv22z4 = (~(vis_r12_o[27] & N71xx4));
assign Ct22z4 = (Uv22z4 & Bw22z4);
assign Bw22z4 = (Iw22z4 & Pw22z4);
assign Pw22z4 = (~(vis_r11_o[27] & Y91xx4));
assign Iw22z4 = (~(vis_r10_o[27] & Ld1xx4));
assign Uv22z4 = (Ww22z4 & Dx22z4);
assign Dx22z4 = (~(vis_r9_o[27] & Ab1xx4));
assign Ww22z4 = (~(vis_r8_o[27] & Sd1xx4));
assign Os22z4 = (Kx22z4 & Rx22z4);
assign Rx22z4 = (Yx22z4 & Fy22z4);
assign Fy22z4 = (My22z4 & Ty22z4);
assign Ty22z4 = (~(vis_r7_o[27] & Jc1xx4));
assign My22z4 = (~(vis_r6_o[27] & T31xx4));
assign Yx22z4 = (Az22z4 & Hz22z4);
assign Hz22z4 = (~(vis_r5_o[27] & U71xx4));
assign Az22z4 = (~(vis_r4_o[27] & R91xx4));
assign Kx22z4 = (Oz22z4 & Vz22z4);
assign Vz22z4 = (C032z4 & J032z4);
assign J032z4 = (~(vis_r3_o[27] & Qc1xx4));
assign C032z4 = (~(vis_r2_o[27] & S61xx4));
assign Oz22z4 = (Q032z4 & X032z4);
assign X032z4 = (~(vis_r1_o[27] & V41xx4));
assign Q032z4 = (~(vis_r0_o[27] & A41xx4));
assign hwdata_o[26] = (~(E132z4 & L132z4));
assign L132z4 = (~(N01xx4 & Zh5wx4));
assign Zh5wx4 = (~(S132z4 & Z132z4));
assign Z132z4 = (G232z4 & N232z4);
assign N232z4 = (U232z4 & B332z4);
assign B332z4 = (I332z4 & P332z4);
assign P332z4 = (~(Gcdvx4 & Ta1xx4));
assign I332z4 = (W332z4 & D432z4);
assign D432z4 = (~(vis_psp_o[8] & Y21xx4));
assign W332z4 = (~(vis_msp_o[8] & C51xx4));
assign U232z4 = (K432z4 & R432z4);
assign R432z4 = (~(vis_r14_o[10] & L61xx4));
assign K432z4 = (~(vis_r12_o[10] & N71xx4));
assign G232z4 = (Y432z4 & F532z4);
assign F532z4 = (M532z4 & T532z4);
assign T532z4 = (~(vis_r11_o[10] & Y91xx4));
assign M532z4 = (~(vis_r10_o[10] & Ld1xx4));
assign Y432z4 = (A632z4 & H632z4);
assign H632z4 = (~(vis_r9_o[10] & Ab1xx4));
assign A632z4 = (~(vis_r8_o[10] & Sd1xx4));
assign S132z4 = (O632z4 & V632z4);
assign V632z4 = (C732z4 & J732z4);
assign J732z4 = (Q732z4 & X732z4);
assign X732z4 = (~(vis_r7_o[10] & Jc1xx4));
assign Q732z4 = (~(vis_r6_o[10] & T31xx4));
assign C732z4 = (E832z4 & L832z4);
assign L832z4 = (~(vis_r5_o[10] & U71xx4));
assign E832z4 = (~(vis_r4_o[10] & R91xx4));
assign O632z4 = (S832z4 & Z832z4);
assign Z832z4 = (G932z4 & N932z4);
assign N932z4 = (~(vis_r3_o[10] & Qc1xx4));
assign G932z4 = (~(vis_r2_o[10] & S61xx4));
assign S832z4 = (U932z4 & Ba32z4);
assign Ba32z4 = (~(vis_r1_o[10] & V41xx4));
assign U932z4 = (~(vis_r0_o[10] & A41xx4));
assign E132z4 = (Ia32z4 & Pa32z4);
assign Pa32z4 = (~(Wq5wx4 & Sh5wx4));
assign Sh5wx4 = (~(Wa32z4 & Db32z4));
assign Db32z4 = (Kb32z4 & Rb32z4);
assign Rb32z4 = (Yb32z4 & Fc32z4);
assign Fc32z4 = (~(E1dvx4 & Ta1xx4));
assign Yb32z4 = (Mc32z4 & Tc32z4);
assign Tc32z4 = (~(vis_psp_o[0] & Y21xx4));
assign Mc32z4 = (~(vis_msp_o[0] & C51xx4));
assign Kb32z4 = (Ad32z4 & Hd32z4);
assign Hd32z4 = (~(vis_r14_o[2] & L61xx4));
assign Ad32z4 = (~(vis_r12_o[2] & N71xx4));
assign Wa32z4 = (Od32z4 & Vd32z4);
assign Vd32z4 = (Ce32z4 & Je32z4);
assign Je32z4 = (~(vis_r9_o[2] & Ab1xx4));
assign Ce32z4 = (Qe32z4 & Xe32z4);
assign Xe32z4 = (~(vis_r11_o[2] & Y91xx4));
assign Qe32z4 = (~(vis_r10_o[2] & Ld1xx4));
assign Od32z4 = (Q1ywx4 & Ef32z4);
assign Ef32z4 = (~(vis_r8_o[2] & Sd1xx4));
assign Q1ywx4 = (Lf32z4 & Sf32z4);
assign Sf32z4 = (Zf32z4 & Gg32z4);
assign Gg32z4 = (Ng32z4 & Ug32z4);
assign Ug32z4 = (~(vis_r2_o[2] & S61xx4));
assign Ng32z4 = (~(vis_r6_o[2] & T31xx4));
assign Zf32z4 = (Bh32z4 & Ih32z4);
assign Ih32z4 = (~(vis_r5_o[2] & U71xx4));
assign Bh32z4 = (~(vis_r4_o[2] & R91xx4));
assign Lf32z4 = (Ph32z4 & Wh32z4);
assign Wh32z4 = (Di32z4 & Ki32z4);
assign Ki32z4 = (~(vis_r1_o[2] & V41xx4));
assign Di32z4 = (~(vis_r0_o[2] & A41xx4));
assign Ph32z4 = (Ri32z4 & Yi32z4);
assign Yi32z4 = (~(vis_r3_o[2] & Qc1xx4));
assign Ri32z4 = (~(vis_r7_o[2] & Jc1xx4));
assign Ia32z4 = (~(Ge1xx4 & Pg8wx4));
assign Pg8wx4 = (!Djzvx4);
assign Djzvx4 = (Fj32z4 & Mj32z4);
assign Mj32z4 = (Tj32z4 & Ak32z4);
assign Ak32z4 = (Hk32z4 & Ok32z4);
assign Ok32z4 = (Vk32z4 & Cl32z4);
assign Cl32z4 = (~(Azdvx4 & Ta1xx4));
assign Vk32z4 = (Jl32z4 & Ql32z4);
assign Ql32z4 = (~(vis_psp_o[24] & Y21xx4));
assign Jl32z4 = (~(vis_msp_o[24] & C51xx4));
assign Hk32z4 = (Xl32z4 & Em32z4);
assign Em32z4 = (~(vis_r14_o[26] & L61xx4));
assign Xl32z4 = (~(vis_r12_o[26] & N71xx4));
assign Tj32z4 = (Lm32z4 & Sm32z4);
assign Sm32z4 = (Zm32z4 & Gn32z4);
assign Gn32z4 = (~(vis_r11_o[26] & Y91xx4));
assign Zm32z4 = (~(vis_r10_o[26] & Ld1xx4));
assign Lm32z4 = (Nn32z4 & Un32z4);
assign Un32z4 = (~(vis_r9_o[26] & Ab1xx4));
assign Nn32z4 = (~(vis_r8_o[26] & Sd1xx4));
assign Fj32z4 = (Bo32z4 & Io32z4);
assign Io32z4 = (Po32z4 & Wo32z4);
assign Wo32z4 = (Dp32z4 & Kp32z4);
assign Kp32z4 = (~(vis_r7_o[26] & Jc1xx4));
assign Dp32z4 = (~(vis_r6_o[26] & T31xx4));
assign Po32z4 = (Rp32z4 & Yp32z4);
assign Yp32z4 = (~(vis_r5_o[26] & U71xx4));
assign Rp32z4 = (~(vis_r4_o[26] & R91xx4));
assign Bo32z4 = (Fq32z4 & Mq32z4);
assign Mq32z4 = (Tq32z4 & Ar32z4);
assign Ar32z4 = (~(vis_r3_o[26] & Qc1xx4));
assign Tq32z4 = (~(vis_r2_o[26] & S61xx4));
assign Fq32z4 = (Hr32z4 & Or32z4);
assign Or32z4 = (~(vis_r1_o[26] & V41xx4));
assign Hr32z4 = (~(vis_r0_o[26] & A41xx4));
assign hwdata_o[25] = (~(Vr32z4 & Cs32z4));
assign Cs32z4 = (~(N01xx4 & Vf5wx4));
assign Vf5wx4 = (~(Js32z4 & Qs32z4));
assign Qs32z4 = (Xs32z4 & Et32z4);
assign Et32z4 = (Lt32z4 & St32z4);
assign St32z4 = (Zt32z4 & Gu32z4);
assign Gu32z4 = (~(Wadvx4 & Ta1xx4));
assign Zt32z4 = (Nu32z4 & Uu32z4);
assign Uu32z4 = (~(vis_psp_o[7] & Y21xx4));
assign Nu32z4 = (~(vis_msp_o[7] & C51xx4));
assign Lt32z4 = (Bv32z4 & Iv32z4);
assign Iv32z4 = (~(vis_r14_o[9] & L61xx4));
assign Bv32z4 = (~(vis_r12_o[9] & N71xx4));
assign Xs32z4 = (Pv32z4 & Wv32z4);
assign Wv32z4 = (Dw32z4 & Kw32z4);
assign Kw32z4 = (~(vis_r11_o[9] & Y91xx4));
assign Dw32z4 = (~(vis_r10_o[9] & Ld1xx4));
assign Pv32z4 = (Rw32z4 & Yw32z4);
assign Yw32z4 = (~(vis_r9_o[9] & Ab1xx4));
assign Rw32z4 = (~(vis_r8_o[9] & Sd1xx4));
assign Js32z4 = (Fx32z4 & Mx32z4);
assign Mx32z4 = (Tx32z4 & Ay32z4);
assign Ay32z4 = (Hy32z4 & Oy32z4);
assign Oy32z4 = (~(vis_r7_o[9] & Jc1xx4));
assign Hy32z4 = (~(vis_r6_o[9] & T31xx4));
assign Tx32z4 = (Vy32z4 & Cz32z4);
assign Cz32z4 = (~(vis_r5_o[9] & U71xx4));
assign Vy32z4 = (~(vis_r4_o[9] & R91xx4));
assign Fx32z4 = (Jz32z4 & Qz32z4);
assign Qz32z4 = (Xz32z4 & E042z4);
assign E042z4 = (~(vis_r3_o[9] & Qc1xx4));
assign Xz32z4 = (~(vis_r2_o[9] & S61xx4));
assign Jz32z4 = (L042z4 & S042z4);
assign S042z4 = (~(vis_r1_o[9] & V41xx4));
assign L042z4 = (~(vis_r0_o[9] & A41xx4));
assign Vr32z4 = (Z042z4 & G142z4);
assign G142z4 = (~(Wq5wx4 & Htyvx4));
assign Htyvx4 = (~(N142z4 & U142z4));
assign U142z4 = (B242z4 & I242z4);
assign I242z4 = (P242z4 & W242z4);
assign W242z4 = (~(Uzcvx4 & Ta1xx4));
assign P242z4 = (~(vis_r14_o[1] & L61xx4));
assign B242z4 = (D342z4 & K342z4);
assign K342z4 = (~(vis_r12_o[1] & N71xx4));
assign D342z4 = (~(vis_r11_o[1] & Y91xx4));
assign N142z4 = (R342z4 & Y342z4);
assign Y342z4 = (F442z4 & M442z4);
assign M442z4 = (~(vis_r10_o[1] & Ld1xx4));
assign F442z4 = (~(vis_r9_o[1] & Ab1xx4));
assign R342z4 = (V7ywx4 & T442z4);
assign T442z4 = (~(vis_r8_o[1] & Sd1xx4));
assign V7ywx4 = (A542z4 & H542z4);
assign H542z4 = (O542z4 & V542z4);
assign V542z4 = (C642z4 & J642z4);
assign J642z4 = (~(vis_r7_o[1] & Jc1xx4));
assign C642z4 = (~(vis_r6_o[1] & T31xx4));
assign O542z4 = (Q642z4 & X642z4);
assign X642z4 = (~(vis_r5_o[1] & U71xx4));
assign Q642z4 = (~(vis_r4_o[1] & R91xx4));
assign A542z4 = (E742z4 & L742z4);
assign L742z4 = (S742z4 & Z742z4);
assign Z742z4 = (~(vis_r3_o[1] & Qc1xx4));
assign S742z4 = (~(vis_r2_o[1] & S61xx4));
assign E742z4 = (G842z4 & N842z4);
assign N842z4 = (~(vis_r1_o[1] & V41xx4));
assign G842z4 = (~(vis_r0_o[1] & A41xx4));
assign Z042z4 = (~(Ge1xx4 & Ig8wx4));
assign Ig8wx4 = (!Kqzvx4);
assign Kqzvx4 = (U842z4 & B942z4);
assign B942z4 = (I942z4 & P942z4);
assign P942z4 = (W942z4 & Da42z4);
assign Da42z4 = (Ka42z4 & Ra42z4);
assign Ra42z4 = (~(Pxdvx4 & Ta1xx4));
assign Ka42z4 = (Ya42z4 & Fb42z4);
assign Fb42z4 = (~(vis_psp_o[23] & Y21xx4));
assign Ya42z4 = (~(vis_msp_o[23] & C51xx4));
assign W942z4 = (Mb42z4 & Tb42z4);
assign Tb42z4 = (~(vis_r14_o[25] & L61xx4));
assign Mb42z4 = (~(vis_r12_o[25] & N71xx4));
assign I942z4 = (Ac42z4 & Hc42z4);
assign Hc42z4 = (Oc42z4 & Vc42z4);
assign Vc42z4 = (~(vis_r11_o[25] & Y91xx4));
assign Oc42z4 = (~(vis_r10_o[25] & Ld1xx4));
assign Ac42z4 = (Cd42z4 & Jd42z4);
assign Jd42z4 = (~(vis_r9_o[25] & Ab1xx4));
assign Cd42z4 = (~(vis_r8_o[25] & Sd1xx4));
assign U842z4 = (Qd42z4 & Xd42z4);
assign Xd42z4 = (Ee42z4 & Le42z4);
assign Le42z4 = (Se42z4 & Ze42z4);
assign Ze42z4 = (~(vis_r7_o[25] & Jc1xx4));
assign Se42z4 = (~(vis_r6_o[25] & T31xx4));
assign Ee42z4 = (Gf42z4 & Nf42z4);
assign Nf42z4 = (~(vis_r5_o[25] & U71xx4));
assign Gf42z4 = (~(vis_r4_o[25] & R91xx4));
assign Qd42z4 = (Uf42z4 & Bg42z4);
assign Bg42z4 = (Ig42z4 & Pg42z4);
assign Pg42z4 = (~(vis_r3_o[25] & Qc1xx4));
assign Ig42z4 = (~(vis_r2_o[25] & S61xx4));
assign Uf42z4 = (Wg42z4 & Dh42z4);
assign Dh42z4 = (~(vis_r1_o[25] & V41xx4));
assign Wg42z4 = (~(vis_r0_o[25] & A41xx4));
assign hwdata_o[24] = (~(Kh42z4 & Rh42z4));
assign Rh42z4 = (~(N01xx4 & Rd5wx4));
assign Rd5wx4 = (!P12wx4);
assign P12wx4 = (Yh42z4 & Fi42z4);
assign Fi42z4 = (Mi42z4 & Ti42z4);
assign Ti42z4 = (Aj42z4 & Hj42z4);
assign Hj42z4 = (Oj42z4 & Vj42z4);
assign Vj42z4 = (~(vis_psp_o[6] & Y21xx4));
assign Oj42z4 = (Ck42z4 & Jk42z4);
assign Jk42z4 = (~(vis_r6_o[8] & T31xx4));
assign Ck42z4 = (~(vis_r0_o[8] & A41xx4));
assign Aj42z4 = (Qk42z4 & Xk42z4);
assign Xk42z4 = (~(vis_r1_o[8] & V41xx4));
assign Qk42z4 = (~(vis_msp_o[6] & C51xx4));
assign Mi42z4 = (El42z4 & Ll42z4);
assign Ll42z4 = (Sl42z4 & Zl42z4);
assign Zl42z4 = (~(vis_r14_o[8] & L61xx4));
assign Sl42z4 = (~(vis_r2_o[8] & S61xx4));
assign El42z4 = (Gm42z4 & Nm42z4);
assign Nm42z4 = (~(vis_r12_o[8] & N71xx4));
assign Gm42z4 = (~(vis_r5_o[8] & U71xx4));
assign Yh42z4 = (Um42z4 & Bn42z4);
assign Bn42z4 = (In42z4 & Pn42z4);
assign Pn42z4 = (Wn42z4 & Do42z4);
assign Do42z4 = (~(vis_r4_o[8] & R91xx4));
assign Wn42z4 = (~(vis_r11_o[8] & Y91xx4));
assign In42z4 = (Ko42z4 & Ro42z4);
assign Ro42z4 = (~(M9dvx4 & Ta1xx4));
assign Ko42z4 = (~(vis_r9_o[8] & Ab1xx4));
assign Um42z4 = (Yo42z4 & Fp42z4);
assign Fp42z4 = (Mp42z4 & Tp42z4);
assign Tp42z4 = (~(vis_r7_o[8] & Jc1xx4));
assign Mp42z4 = (~(vis_r3_o[8] & Qc1xx4));
assign Yo42z4 = (Aq42z4 & Hq42z4);
assign Hq42z4 = (~(vis_r10_o[8] & Ld1xx4));
assign Aq42z4 = (~(vis_r8_o[8] & Sd1xx4));
assign N01xx4 = (Oq42z4 & Pp8vx4);
assign Kh42z4 = (Vq42z4 & Cr42z4);
assign Cr42z4 = (Yd5wx4 | Zhyvx4);
assign Yd5wx4 = (!Wq5wx4);
assign Wq5wx4 = (Jr42z4 & Qr42z4);
assign Jr42z4 = (~(C5vvx4 | Oq42z4));
assign Vq42z4 = (~(Ge1xx4 & Eacwx4));
assign Eacwx4 = (~(Xr42z4 & Es42z4));
assign Es42z4 = (Ls42z4 & Ss42z4);
assign Ss42z4 = (Zs42z4 & Gt42z4);
assign Gt42z4 = (Nt42z4 & Ut42z4);
assign Ut42z4 = (~(Ewdvx4 & Ta1xx4));
assign Nt42z4 = (Bu42z4 & Iu42z4);
assign Iu42z4 = (~(vis_psp_o[22] & Y21xx4));
assign Bu42z4 = (~(vis_msp_o[22] & C51xx4));
assign Zs42z4 = (Pu42z4 & Wu42z4);
assign Wu42z4 = (~(vis_r14_o[24] & L61xx4));
assign Pu42z4 = (~(vis_r12_o[24] & N71xx4));
assign Ls42z4 = (Dv42z4 & Kv42z4);
assign Kv42z4 = (Rv42z4 & Yv42z4);
assign Yv42z4 = (~(vis_r11_o[24] & Y91xx4));
assign Rv42z4 = (~(vis_r10_o[24] & Ld1xx4));
assign Dv42z4 = (Fw42z4 & Mw42z4);
assign Mw42z4 = (~(vis_r9_o[24] & Ab1xx4));
assign Fw42z4 = (~(vis_r8_o[24] & Sd1xx4));
assign Xr42z4 = (Tw42z4 & Ax42z4);
assign Ax42z4 = (Hx42z4 & Ox42z4);
assign Ox42z4 = (Vx42z4 & Cy42z4);
assign Cy42z4 = (~(vis_r7_o[24] & Jc1xx4));
assign Vx42z4 = (~(vis_r6_o[24] & T31xx4));
assign Hx42z4 = (Jy42z4 & Qy42z4);
assign Qy42z4 = (~(vis_r5_o[24] & U71xx4));
assign Jy42z4 = (~(vis_r4_o[24] & R91xx4));
assign Tw42z4 = (Xy42z4 & Ez42z4);
assign Ez42z4 = (Lz42z4 & Sz42z4);
assign Sz42z4 = (~(vis_r3_o[24] & Qc1xx4));
assign Lz42z4 = (~(vis_r2_o[24] & S61xx4));
assign Xy42z4 = (Zz42z4 & G052z4);
assign G052z4 = (~(vis_r1_o[24] & V41xx4));
assign Zz42z4 = (~(vis_r0_o[24] & A41xx4));
assign hwdata_o[23] = (Ge1xx4 ? R6cwx4 : Ht5wx4);
assign Ge1xx4 = (Pp8vx4 & N052z4);
assign N052z4 = (!Qr42z4);
assign R6cwx4 = (~(U052z4 & B152z4));
assign B152z4 = (I152z4 & P152z4);
assign P152z4 = (W152z4 & D252z4);
assign D252z4 = (K252z4 & R252z4);
assign R252z4 = (~(Tudvx4 & Ta1xx4));
assign K252z4 = (Y252z4 & F352z4);
assign F352z4 = (~(vis_psp_o[21] & Y21xx4));
assign Y252z4 = (~(vis_msp_o[21] & C51xx4));
assign W152z4 = (M352z4 & T352z4);
assign T352z4 = (~(vis_r14_o[23] & L61xx4));
assign M352z4 = (~(vis_r12_o[23] & N71xx4));
assign I152z4 = (A452z4 & H452z4);
assign H452z4 = (O452z4 & V452z4);
assign V452z4 = (~(vis_r11_o[23] & Y91xx4));
assign O452z4 = (~(vis_r10_o[23] & Ld1xx4));
assign A452z4 = (C552z4 & J552z4);
assign J552z4 = (~(vis_r9_o[23] & Ab1xx4));
assign C552z4 = (~(vis_r8_o[23] & Sd1xx4));
assign U052z4 = (Q552z4 & X552z4);
assign X552z4 = (E652z4 & L652z4);
assign L652z4 = (S652z4 & Z652z4);
assign Z652z4 = (~(vis_r7_o[23] & Jc1xx4));
assign S652z4 = (~(vis_r6_o[23] & T31xx4));
assign E652z4 = (G752z4 & N752z4);
assign N752z4 = (~(vis_r5_o[23] & U71xx4));
assign G752z4 = (~(vis_r4_o[23] & R91xx4));
assign Q552z4 = (U752z4 & B852z4);
assign B852z4 = (I852z4 & P852z4);
assign P852z4 = (~(vis_r3_o[23] & Qc1xx4));
assign I852z4 = (~(vis_r2_o[23] & S61xx4));
assign U752z4 = (W852z4 & D952z4);
assign D952z4 = (~(vis_r1_o[23] & V41xx4));
assign W852z4 = (~(vis_r0_o[23] & A41xx4));
assign Ht5wx4 = (~(K952z4 & R952z4));
assign R952z4 = (Y952z4 & Fa52z4);
assign Fa52z4 = (Ma52z4 & Ta52z4);
assign Ta52z4 = (~(C8dvx4 & Ta1xx4));
assign Ma52z4 = (Ab52z4 & Hb52z4);
assign Hb52z4 = (~(vis_psp_o[5] & Y21xx4));
assign Y21xx4 = (Ob52z4 & O7evx4);
assign Ob52z4 = (~(Vb52z4 | Cc52z4));
assign Ab52z4 = (~(vis_msp_o[5] & C51xx4));
assign C51xx4 = (Jc52z4 & Qc52z4);
assign Jc52z4 = (~(Cc52z4 | O7evx4));
assign Y952z4 = (Xc52z4 & Ed52z4);
assign Ed52z4 = (~(vis_r14_o[7] & L61xx4));
assign Xc52z4 = (~(vis_r12_o[7] & N71xx4));
assign K952z4 = (Ld52z4 & Sd52z4);
assign Sd52z4 = (Zd52z4 & Ge52z4);
assign Ge52z4 = (~(vis_r9_o[7] & Ab1xx4));
assign Zd52z4 = (Ne52z4 & Ue52z4);
assign Ue52z4 = (~(vis_r11_o[7] & Y91xx4));
assign Ne52z4 = (~(vis_r10_o[7] & Ld1xx4));
assign Ld52z4 = (Xowwx4 & Bf52z4);
assign Bf52z4 = (~(vis_r8_o[7] & Sd1xx4));
assign Xowwx4 = (If52z4 & Pf52z4);
assign Pf52z4 = (Wf52z4 & Dg52z4);
assign Dg52z4 = (Kg52z4 & Rg52z4);
assign Rg52z4 = (~(vis_r0_o[7] & A41xx4));
assign Kg52z4 = (~(vis_r2_o[7] & S61xx4));
assign Wf52z4 = (Yg52z4 & Fh52z4);
assign Fh52z4 = (~(vis_r5_o[7] & U71xx4));
assign Yg52z4 = (~(vis_r4_o[7] & R91xx4));
assign If52z4 = (Mh52z4 & Th52z4);
assign Th52z4 = (Ai52z4 & Hi52z4);
assign Hi52z4 = (~(vis_r7_o[7] & Jc1xx4));
assign Ai52z4 = (~(vis_r3_o[7] & Qc1xx4));
assign Mh52z4 = (Oi52z4 & Vi52z4);
assign Vi52z4 = (~(vis_r1_o[7] & V41xx4));
assign Oi52z4 = (~(vis_r6_o[7] & T31xx4));
assign hwdata_o[0] = (~(C5vvx4 | Zhyvx4));
assign Zhyvx4 = (Cj52z4 & Jj52z4);
assign Jj52z4 = (Qj52z4 & Xj52z4);
assign Xj52z4 = (Ek52z4 & Lk52z4);
assign Lk52z4 = (~(vis_r10_o[0] & Ld1xx4));
assign Ld1xx4 = (~(Sk52z4 | Zk52z4));
assign Ek52z4 = (~(Kycvx4 & Ta1xx4));
assign Ta1xx4 = (~(Gl52z4 | Cc52z4));
assign Qj52z4 = (Nl52z4 & Ul52z4);
assign Ul52z4 = (~(vis_r12_o[0] & N71xx4));
assign N71xx4 = (~(Bm52z4 | Cc52z4));
assign Nl52z4 = (~(vis_r11_o[0] & Y91xx4));
assign Y91xx4 = (~(Sk52z4 | Gl52z4));
assign Cj52z4 = (Im52z4 & Pm52z4);
assign Pm52z4 = (Wm52z4 & Dn52z4);
assign Dn52z4 = (~(vis_r8_o[0] & Sd1xx4));
assign Sd1xx4 = (~(Sk52z4 | Bm52z4));
assign Wm52z4 = (~(vis_r9_o[0] & Ab1xx4));
assign Ab1xx4 = (~(Sk52z4 | Vb52z4));
assign Sk52z4 = (~(Vu8vx4 & Kn52z4));
assign Im52z4 = (Q8ywx4 & Rn52z4);
assign Rn52z4 = (~(vis_r14_o[0] & L61xx4));
assign L61xx4 = (~(Zk52z4 | Cc52z4));
assign Cc52z4 = (~(Vu8vx4 & Nt8vx4));
assign Q8ywx4 = (Yn52z4 & Fo52z4);
assign Fo52z4 = (Mo52z4 & To52z4);
assign To52z4 = (Ap52z4 & Hp52z4);
assign Hp52z4 = (~(vis_r2_o[0] & S61xx4));
assign S61xx4 = (~(Op52z4 | Zk52z4));
assign Ap52z4 = (~(vis_r6_o[0] & T31xx4));
assign T31xx4 = (~(Vp52z4 | Zk52z4));
assign Zk52z4 = (~(Fs8vx4 & Cq52z4));
assign Mo52z4 = (Jq52z4 & Qq52z4);
assign Qq52z4 = (~(vis_r5_o[0] & U71xx4));
assign U71xx4 = (~(Vp52z4 | Vb52z4));
assign Jq52z4 = (~(vis_r4_o[0] & R91xx4));
assign R91xx4 = (~(Vp52z4 | Bm52z4));
assign Yn52z4 = (Xq52z4 & Er52z4);
assign Er52z4 = (Lr52z4 & Sr52z4);
assign Sr52z4 = (~(vis_r1_o[0] & V41xx4));
assign V41xx4 = (~(Op52z4 | Vb52z4));
assign Vb52z4 = (!Qc52z4);
assign Qc52z4 = (Xq8vx4 & Zr52z4);
assign Lr52z4 = (~(vis_r0_o[0] & A41xx4));
assign A41xx4 = (~(Op52z4 | Bm52z4));
assign Bm52z4 = (~(Cq52z4 & Zr52z4));
assign Zr52z4 = (!Fs8vx4);
assign Cq52z4 = (!Xq8vx4);
assign Xq52z4 = (Gs52z4 & Ns52z4);
assign Ns52z4 = (~(vis_r3_o[0] & Qc1xx4));
assign Qc1xx4 = (~(Op52z4 | Gl52z4));
assign Op52z4 = (Nt8vx4 | Vu8vx4);
assign Gs52z4 = (~(vis_r7_o[0] & Jc1xx4));
assign Jc1xx4 = (~(Vp52z4 | Gl52z4));
assign Gl52z4 = (~(Fs8vx4 & Xq8vx4));
assign Vp52z4 = (Kn52z4 | Vu8vx4);
assign Kn52z4 = (!Nt8vx4);
assign C5vvx4 = (!Pp8vx4);
assign htrans_o[1] = (Us52z4 & Xmywx4);
assign Xmywx4 = (E7mwx4 | hprot_o[3]);
assign Us52z4 = (~(Bt52z4 & E7mwx4));
assign E7mwx4 = (It52z4 | hprot_o[0]);
assign hprot_o[0] = (~(Pt52z4 & Wt52z4));
assign Wt52z4 = (Du52z4 & Ku52z4);
assign Ku52z4 = (Ru52z4 & Z0mwx4);
assign Z0mwx4 = (~(Yu52z4 | Fv52z4));
assign Fv52z4 = (Mv52z4 & Ibdwx4);
assign Ibdwx4 = (~(U9gvx4 | Whgvx4));
assign Mv52z4 = (B73wx4 & S4xvx4);
assign Yu52z4 = (Tv52z4 & Xhqvx4);
assign Tv52z4 = (~(S87wx4 | F3ovx4));
assign Du52z4 = (Aw52z4 & Mrkwx4);
assign Mrkwx4 = (~(Hw52z4 & Huqvx4));
assign Hw52z4 = (Kzxvx4 & Hgxvx4);
assign Aw52z4 = (A76wx4 & Yy5wx4);
assign Yy5wx4 = (~(Ow52z4 & O76wx4));
assign Ow52z4 = (~(J43wx4 | Vdgvx4));
assign A76wx4 = (~(Clewx4 & R5dwx4));
assign Pt52z4 = (Vw52z4 & Cx52z4);
assign Cx52z4 = (Jx52z4 & Qx52z4);
assign Qx52z4 = (~(Xx52z4 & Ey52z4));
assign Ey52z4 = (~(Rexvx4 | Mj8vx4));
assign Xx52z4 = (~(Njxvx4 | Us2wx4));
assign Njxvx4 = (!Liqvx4);
assign Liqvx4 = (~(Hq1wx4 | Zrvvx4));
assign Jx52z4 = (Ly52z4 & Sy52z4);
assign Sy52z4 = (~(Zy52z4 & Ilhwx4));
assign Ilhwx4 = (~(S4xvx4 | Dmgvx4));
assign Zy52z4 = (~(Pxyvx4 | Nggvx4));
assign Ly52z4 = (~(Zmewx4 & O9qvx4));
assign Vw52z4 = (Gz52z4 & Ol6wx4);
assign Gz52z4 = (Nz52z4 & Uz52z4);
assign Uz52z4 = (~(T1xvx4 & Cihwx4));
assign Cihwx4 = (~(Q5gvx4 | Mcgvx4));
assign Nz52z4 = (~(B062z4 & Clewx4));
assign B062z4 = (~(F3ovx4 | Vdgvx4));
assign Bt52z4 = (~(I062z4 & P062z4));
assign P062z4 = (~(W062z4 | W6qvx4));
assign W6qvx4 = (D162z4 & K162z4);
assign K162z4 = (~(V3wvx4 & R162z4));
assign R162z4 = (~(Y162z4 & T50wx4));
assign D162z4 = (Y162z4 | Oq42z4);
assign W062z4 = (Trsvx4 | Mrsvx4);
assign I062z4 = (Ppsvx4 & F262z4);
assign F262z4 = (~(Hssvx4 & V2qvx4));
assign Hssvx4 = (M262z4 & haddr_o[31]);
assign M262z4 = (haddr_o[30] & haddr_o[29]);
assign hsize_o[1] = (~(It52z4 & T262z4));
assign T262z4 = (Qr42z4 | Mrsvx4);
assign hsize_o[0] = (A362z4 & Oq42z4);
assign A362z4 = (It52z4 & D7qvx4);
assign hprot_o[3] = (~(hprot_o[2] & H362z4));
assign H362z4 = (~(O362z4 & V362z4));
assign V362z4 = (~(C462z4 & J462z4));
assign J462z4 = (Ovpvx4 | Ykh2z4[30]);
assign Ovpvx4 = (!haddr_o[29]);
assign C462z4 = (~(Q462z4 | X462z4));
assign hprot_o[2] = (haddr_o[30] | haddr_o[29]);
assign haddr_o[29] = (E562z4 | Q462z4);
assign Q462z4 = (Gzvvx4 & Xrnvx4);
assign Xrnvx4 = (~(L562z4 & S562z4));
assign S562z4 = (~(W1evx4 & Jj9wx4));
assign L562z4 = (Z562z4 & G662z4);
assign G662z4 = (~(Vb9wx4 & N662z4));
assign N662z4 = (~(U662z4 & B762z4));
assign B762z4 = (I762z4 & P762z4);
assign P762z4 = (W762z4 & D862z4);
assign D862z4 = (~(vis_r14_o[29] & Zd9wx4));
assign W762z4 = (K862z4 & R862z4);
assign R862z4 = (~(vis_psp_o[27] & Ue9wx4));
assign K862z4 = (~(vis_msp_o[27] & Bf9wx4));
assign I762z4 = (Y862z4 & F962z4);
assign F962z4 = (~(vis_r12_o[29] & Wf9wx4));
assign Y862z4 = (~(vis_r11_o[29] & Dg9wx4));
assign U662z4 = (M962z4 & T962z4);
assign T962z4 = (Aa62z4 & Ha62z4);
assign Ha62z4 = (~(vis_r10_o[29] & Mh9wx4));
assign Aa62z4 = (~(vis_r9_o[29] & Th9wx4));
assign M962z4 = (Eruwx4 & Oa62z4);
assign Oa62z4 = (~(vis_r8_o[29] & Oi9wx4));
assign Z562z4 = (~(H3evx4 & Qj9wx4));
assign E562z4 = (X462z4 | Va62z4);
assign Va62z4 = (Ykh2z4[28] & Mrsvx4);
assign X462z4 = (Dmh2z4[29] & K1wvx4);
assign haddr_o[30] = (~(Cb62z4 & Jb62z4));
assign Jb62z4 = (~(Gzvvx4 & Hqnvx4));
assign Hqnvx4 = (!Q8zvx4);
assign Q8zvx4 = (Qb62z4 & Xb62z4);
assign Xb62z4 = (~(Vb9wx4 & Ec62z4));
assign Ec62z4 = (~(Lc62z4 & Sc62z4));
assign Sc62z4 = (Zc62z4 & Gd62z4);
assign Gd62z4 = (Nd62z4 & Ud62z4);
assign Ud62z4 = (~(vis_r14_o[30] & Zd9wx4));
assign Nd62z4 = (Be62z4 & Ie62z4);
assign Ie62z4 = (~(vis_psp_o[28] & Ue9wx4));
assign Be62z4 = (~(vis_msp_o[28] & Bf9wx4));
assign Zc62z4 = (Pe62z4 & We62z4);
assign We62z4 = (~(vis_r12_o[30] & Wf9wx4));
assign Pe62z4 = (~(vis_r11_o[30] & Dg9wx4));
assign Lc62z4 = (Df62z4 & Kf62z4);
assign Kf62z4 = (Rf62z4 & Yf62z4);
assign Yf62z4 = (~(vis_r10_o[30] & Mh9wx4));
assign Rf62z4 = (~(vis_r9_o[30] & Th9wx4));
assign Df62z4 = (Saqwx4 & Fg62z4);
assign Fg62z4 = (~(vis_r8_o[30] & Oi9wx4));
assign Qb62z4 = (Mg62z4 & Tg62z4);
assign Tg62z4 = (~(H3evx4 & Jj9wx4));
assign Mg62z4 = (~(S4evx4 & Qj9wx4));
assign Cb62z4 = (Ah62z4 & Hh62z4);
assign Hh62z4 = (~(Ykh2z4[29] & Mrsvx4));
assign Ah62z4 = (~(Dmh2z4[30] & K1wvx4));
assign haddr_o[7] = (!S4qvx4);
assign S4qvx4 = (Oh62z4 & Vh62z4);
assign Vh62z4 = (~(Ykh2z4[6] & Mrsvx4));
assign Oh62z4 = (Ci62z4 & Ji62z4);
assign Ji62z4 = (~(Gzvvx4 & Yonvx4));
assign Yonvx4 = (~(Qi62z4 & Xi62z4));
assign Xi62z4 = (~(S6dvx4 & Jj9wx4));
assign Qi62z4 = (Ej62z4 & Lj62z4);
assign Lj62z4 = (~(Vb9wx4 & Sj62z4));
assign Sj62z4 = (~(Zj62z4 & Gk62z4));
assign Gk62z4 = (Nk62z4 & Uk62z4);
assign Uk62z4 = (Bl62z4 & Il62z4);
assign Il62z4 = (~(Zd9wx4 & vis_r14_o[7]));
assign Bl62z4 = (Pl62z4 & Wl62z4);
assign Wl62z4 = (~(Ue9wx4 & vis_psp_o[5]));
assign Pl62z4 = (~(Bf9wx4 & vis_msp_o[5]));
assign Nk62z4 = (Dm62z4 & Km62z4);
assign Km62z4 = (~(Wf9wx4 & vis_r12_o[7]));
assign Dm62z4 = (~(Dg9wx4 & vis_r11_o[7]));
assign Zj62z4 = (Rm62z4 & Ym62z4);
assign Ym62z4 = (Fn62z4 & Mn62z4);
assign Mn62z4 = (~(Mh9wx4 & vis_r10_o[7]));
assign Fn62z4 = (~(Th9wx4 & vis_r9_o[7]));
assign Rm62z4 = (Bywwx4 & Tn62z4);
assign Tn62z4 = (~(Oi9wx4 & vis_r8_o[7]));
assign Ej62z4 = (~(Qj9wx4 & C8dvx4));
assign Ci62z4 = (~(Dmh2z4[7] & K1wvx4));
assign haddr_o[6] = (!Hszvx4);
assign Hszvx4 = (Ao62z4 & Ho62z4);
assign Ho62z4 = (~(Ykh2z4[5] & Mrsvx4));
assign Ao62z4 = (Oo62z4 & Vo62z4);
assign Vo62z4 = (~(Gzvvx4 & Fpnvx4));
assign Fpnvx4 = (!Euzvx4);
assign Euzvx4 = (Cp62z4 & Jp62z4);
assign Jp62z4 = (~(Vb9wx4 & Qp62z4));
assign Qp62z4 = (~(Xp62z4 & Eq62z4));
assign Eq62z4 = (Lq62z4 & Sq62z4);
assign Sq62z4 = (Zq62z4 & Gr62z4);
assign Gr62z4 = (~(Zd9wx4 & vis_r14_o[6]));
assign Zq62z4 = (Nr62z4 & Ur62z4);
assign Ur62z4 = (~(Ue9wx4 & vis_psp_o[4]));
assign Nr62z4 = (~(Bf9wx4 & vis_msp_o[4]));
assign Lq62z4 = (Bs62z4 & Is62z4);
assign Is62z4 = (~(Wf9wx4 & vis_r12_o[6]));
assign Bs62z4 = (~(Dg9wx4 & vis_r11_o[6]));
assign Xp62z4 = (Ps62z4 & Ws62z4);
assign Ws62z4 = (Dt62z4 & Kt62z4);
assign Kt62z4 = (~(Mh9wx4 & vis_r10_o[6]));
assign Dt62z4 = (~(Th9wx4 & vis_r9_o[6]));
assign Ps62z4 = (Svqwx4 & Rt62z4);
assign Rt62z4 = (~(Oi9wx4 & vis_r8_o[6]));
assign Cp62z4 = (Yt62z4 & Fu62z4);
assign Fu62z4 = (~(I5dvx4 & Jj9wx4));
assign Yt62z4 = (~(Qj9wx4 & S6dvx4));
assign Oo62z4 = (~(Dmh2z4[6] & K1wvx4));
assign haddr_o[5] = (!Rxzvx4);
assign Rxzvx4 = (Mu62z4 & Tu62z4);
assign Tu62z4 = (~(Ykh2z4[4] & Mrsvx4));
assign Mu62z4 = (Av62z4 & Hv62z4);
assign Hv62z4 = (~(Gzvvx4 & Mpnvx4));
assign Mpnvx4 = (~(Ov62z4 & Vv62z4));
assign Vv62z4 = (~(Y3dvx4 & Jj9wx4));
assign Ov62z4 = (Cw62z4 & Jw62z4);
assign Jw62z4 = (~(Vb9wx4 & Qw62z4));
assign Qw62z4 = (~(Xw62z4 & Ex62z4));
assign Ex62z4 = (Lx62z4 & Sx62z4);
assign Sx62z4 = (Zx62z4 & Gy62z4);
assign Gy62z4 = (~(vis_r14_o[5] & Zd9wx4));
assign Zx62z4 = (Ny62z4 & Uy62z4);
assign Uy62z4 = (~(vis_psp_o[3] & Ue9wx4));
assign Ny62z4 = (~(vis_msp_o[3] & Bf9wx4));
assign Lx62z4 = (Bz62z4 & Iz62z4);
assign Iz62z4 = (~(vis_r12_o[5] & Wf9wx4));
assign Bz62z4 = (~(vis_r11_o[5] & Dg9wx4));
assign Xw62z4 = (Pz62z4 & Wz62z4);
assign Wz62z4 = (D072z4 & K072z4);
assign K072z4 = (~(vis_r10_o[5] & Mh9wx4));
assign D072z4 = (~(vis_r9_o[5] & Th9wx4));
assign Pz62z4 = (Qxuwx4 & R072z4);
assign R072z4 = (~(vis_r8_o[5] & Oi9wx4));
assign Cw62z4 = (~(I5dvx4 & Qj9wx4));
assign Av62z4 = (~(Dmh2z4[5] & K1wvx4));
assign haddr_o[4] = (!Yuovx4);
assign Yuovx4 = (Y072z4 & F172z4);
assign F172z4 = (~(Ykh2z4[3] & Mrsvx4));
assign Y072z4 = (M172z4 & T172z4);
assign T172z4 = (~(Gzvvx4 & Tpnvx4));
assign Tpnvx4 = (~(A272z4 & H272z4));
assign H272z4 = (~(O2dvx4 & Jj9wx4));
assign A272z4 = (O272z4 & V272z4);
assign V272z4 = (~(Vb9wx4 & C372z4));
assign C372z4 = (~(J372z4 & Q372z4));
assign Q372z4 = (X372z4 & E472z4);
assign E472z4 = (L472z4 & S472z4);
assign S472z4 = (~(vis_r14_o[4] & Zd9wx4));
assign L472z4 = (Z472z4 & G572z4);
assign G572z4 = (~(vis_psp_o[2] & Ue9wx4));
assign Z472z4 = (~(vis_msp_o[2] & Bf9wx4));
assign X372z4 = (N572z4 & U572z4);
assign U572z4 = (~(vis_r12_o[4] & Wf9wx4));
assign N572z4 = (~(vis_r11_o[4] & Dg9wx4));
assign J372z4 = (B672z4 & I672z4);
assign I672z4 = (P672z4 & W672z4);
assign W672z4 = (~(vis_r10_o[4] & Mh9wx4));
assign P672z4 = (~(vis_r9_o[4] & Th9wx4));
assign B672z4 = (Bdwwx4 & D772z4);
assign D772z4 = (~(vis_r8_o[4] & Oi9wx4));
assign O272z4 = (~(Y3dvx4 & Qj9wx4));
assign M172z4 = (~(Dmh2z4[4] & K1wvx4));
assign haddr_o[31] = (~(O362z4 & K772z4));
assign K772z4 = (~(Ykh2z4[30] & Mrsvx4));
assign O362z4 = (R772z4 & Y772z4);
assign Y772z4 = (~(Gzvvx4 & A67wx4));
assign A67wx4 = (~(F872z4 & M872z4));
assign M872z4 = (~(S4evx4 & Jj9wx4));
assign F872z4 = (T872z4 & A972z4);
assign A972z4 = (~(Vb9wx4 & H972z4));
assign H972z4 = (~(O972z4 & V972z4));
assign V972z4 = (Ca72z4 & Ja72z4);
assign Ja72z4 = (Qa72z4 & Xa72z4);
assign Xa72z4 = (~(Zd9wx4 & vis_r14_o[31]));
assign Qa72z4 = (Eb72z4 & Lb72z4);
assign Lb72z4 = (~(Ue9wx4 & vis_psp_o[29]));
assign Eb72z4 = (~(Bf9wx4 & vis_msp_o[29]));
assign Ca72z4 = (Sb72z4 & Zb72z4);
assign Zb72z4 = (~(Wf9wx4 & vis_r12_o[31]));
assign Sb72z4 = (~(Dg9wx4 & vis_r11_o[31]));
assign O972z4 = (Gc72z4 & Nc72z4);
assign Nc72z4 = (Uc72z4 & Bd72z4);
assign Bd72z4 = (~(Mh9wx4 & vis_r10_o[31]));
assign Uc72z4 = (~(Th9wx4 & vis_r9_o[31]));
assign Gc72z4 = (N3ywx4 & Id72z4);
assign Id72z4 = (~(Oi9wx4 & vis_r8_o[31]));
assign T872z4 = (~(Qj9wx4 & D6evx4));
assign R772z4 = (~(Dmh2z4[31] & K1wvx4));
assign haddr_o[28] = (!V2qvx4);
assign V2qvx4 = (Pd72z4 & Wd72z4);
assign Wd72z4 = (~(Ykh2z4[27] & Mrsvx4));
assign Pd72z4 = (De72z4 & Ke72z4);
assign Ke72z4 = (~(Gzvvx4 & Esnvx4));
assign Esnvx4 = (~(Re72z4 & Ye72z4));
assign Ye72z4 = (~(L0evx4 & Jj9wx4));
assign Re72z4 = (Ff72z4 & Mf72z4);
assign Mf72z4 = (~(Vb9wx4 & Tf72z4));
assign Tf72z4 = (~(Ag72z4 & Hg72z4));
assign Hg72z4 = (Og72z4 & Vg72z4);
assign Vg72z4 = (Ch72z4 & Jh72z4);
assign Jh72z4 = (~(vis_r14_o[28] & Zd9wx4));
assign Ch72z4 = (Qh72z4 & Xh72z4);
assign Xh72z4 = (~(vis_psp_o[26] & Ue9wx4));
assign Qh72z4 = (~(vis_msp_o[26] & Bf9wx4));
assign Og72z4 = (Ei72z4 & Li72z4);
assign Li72z4 = (~(vis_r12_o[28] & Wf9wx4));
assign Ei72z4 = (~(vis_r11_o[28] & Dg9wx4));
assign Ag72z4 = (Si72z4 & Zi72z4);
assign Zi72z4 = (Gj72z4 & Nj72z4);
assign Nj72z4 = (~(vis_r10_o[28] & Mh9wx4));
assign Gj72z4 = (~(vis_r9_o[28] & Th9wx4));
assign Si72z4 = (F8wwx4 & Uj72z4);
assign Uj72z4 = (~(vis_r8_o[28] & Oi9wx4));
assign Ff72z4 = (~(W1evx4 & Qj9wx4));
assign De72z4 = (~(Dmh2z4[28] & K1wvx4));
assign haddr_o[27] = (!Vezvx4);
assign Vezvx4 = (Bk72z4 & Ik72z4);
assign Ik72z4 = (~(Ykh2z4[26] & Mrsvx4));
assign Bk72z4 = (Pk72z4 & Wk72z4);
assign Wk72z4 = (~(Gzvvx4 & Lsnvx4));
assign Lsnvx4 = (~(Dl72z4 & Kl72z4));
assign Kl72z4 = (~(Azdvx4 & Jj9wx4));
assign Dl72z4 = (Rl72z4 & Yl72z4);
assign Yl72z4 = (~(Vb9wx4 & Fm72z4));
assign Fm72z4 = (~(Mm72z4 & Tm72z4));
assign Tm72z4 = (An72z4 & Hn72z4);
assign Hn72z4 = (On72z4 & Vn72z4);
assign Vn72z4 = (~(vis_r14_o[27] & Zd9wx4));
assign On72z4 = (Co72z4 & Jo72z4);
assign Jo72z4 = (~(vis_psp_o[25] & Ue9wx4));
assign Co72z4 = (~(vis_msp_o[25] & Bf9wx4));
assign An72z4 = (Qo72z4 & Xo72z4);
assign Xo72z4 = (~(vis_r12_o[27] & Wf9wx4));
assign Qo72z4 = (~(vis_r11_o[27] & Dg9wx4));
assign Mm72z4 = (Ep72z4 & Lp72z4);
assign Lp72z4 = (Sp72z4 & Zp72z4);
assign Zp72z4 = (~(vis_r10_o[27] & Mh9wx4));
assign Sp72z4 = (~(vis_r9_o[27] & Th9wx4));
assign Ep72z4 = (Fexwx4 & Gq72z4);
assign Gq72z4 = (~(vis_r8_o[27] & Oi9wx4));
assign Rl72z4 = (~(L0evx4 & Qj9wx4));
assign Pk72z4 = (~(Dmh2z4[27] & K1wvx4));
assign haddr_o[26] = (!Nhzvx4);
assign Nhzvx4 = (Nq72z4 & Uq72z4);
assign Uq72z4 = (~(Ykh2z4[25] & Mrsvx4));
assign Nq72z4 = (Br72z4 & Ir72z4);
assign Ir72z4 = (~(Gzvvx4 & Ssnvx4));
assign Ssnvx4 = (!Hlzvx4);
assign Hlzvx4 = (Pr72z4 & Wr72z4);
assign Wr72z4 = (~(Vb9wx4 & Ds72z4));
assign Ds72z4 = (~(Ks72z4 & Rs72z4));
assign Rs72z4 = (Ys72z4 & Ft72z4);
assign Ft72z4 = (Mt72z4 & Tt72z4);
assign Tt72z4 = (~(Zd9wx4 & vis_r14_o[26]));
assign Mt72z4 = (Au72z4 & Hu72z4);
assign Hu72z4 = (~(Ue9wx4 & vis_psp_o[24]));
assign Au72z4 = (~(Bf9wx4 & vis_msp_o[24]));
assign Ys72z4 = (Ou72z4 & Vu72z4);
assign Vu72z4 = (~(Wf9wx4 & vis_r12_o[26]));
assign Ou72z4 = (~(Dg9wx4 & vis_r11_o[26]));
assign Ks72z4 = (Cv72z4 & Jv72z4);
assign Jv72z4 = (Qv72z4 & Xv72z4);
assign Xv72z4 = (~(Mh9wx4 & vis_r10_o[26]));
assign Qv72z4 = (~(Th9wx4 & vis_r9_o[26]));
assign Cv72z4 = (Feqwx4 & Ew72z4);
assign Ew72z4 = (~(Oi9wx4 & vis_r8_o[26]));
assign Pr72z4 = (Lw72z4 & Sw72z4);
assign Sw72z4 = (~(Pxdvx4 & Jj9wx4));
assign Lw72z4 = (~(Qj9wx4 & Azdvx4));
assign Br72z4 = (~(Dmh2z4[26] & K1wvx4));
assign haddr_o[25] = (!Rnovx4);
assign Rnovx4 = (Zw72z4 & Gx72z4);
assign Gx72z4 = (~(Ykh2z4[24] & Mrsvx4));
assign Zw72z4 = (Nx72z4 & Ux72z4);
assign Ux72z4 = (~(Gzvvx4 & Zsnvx4));
assign Zsnvx4 = (!Nozvx4);
assign Nozvx4 = (By72z4 & Iy72z4);
assign Iy72z4 = (~(Vb9wx4 & Py72z4));
assign Py72z4 = (~(Wy72z4 & Dz72z4));
assign Dz72z4 = (Kz72z4 & Rz72z4);
assign Rz72z4 = (Yz72z4 & F082z4);
assign F082z4 = (~(Zd9wx4 & vis_r14_o[25]));
assign Yz72z4 = (M082z4 & T082z4);
assign T082z4 = (~(Ue9wx4 & vis_psp_o[23]));
assign M082z4 = (~(Bf9wx4 & vis_msp_o[23]));
assign Kz72z4 = (A182z4 & H182z4);
assign H182z4 = (~(Wf9wx4 & vis_r12_o[25]));
assign A182z4 = (~(Dg9wx4 & vis_r11_o[25]));
assign Wy72z4 = (O182z4 & V182z4);
assign V182z4 = (C282z4 & J282z4);
assign J282z4 = (~(Mh9wx4 & vis_r10_o[25]));
assign C282z4 = (~(Th9wx4 & vis_r9_o[25]));
assign O182z4 = (U7uwx4 & Q282z4);
assign Q282z4 = (~(Oi9wx4 & vis_r8_o[25]));
assign By72z4 = (X282z4 & E382z4);
assign E382z4 = (~(Ewdvx4 & Jj9wx4));
assign X282z4 = (~(Qj9wx4 & Pxdvx4));
assign Nx72z4 = (~(Dmh2z4[25] & K1wvx4));
assign haddr_o[24] = (!Y1pvx4);
assign Y1pvx4 = (L382z4 & S382z4);
assign S382z4 = (~(Ykh2z4[23] & Mrsvx4));
assign L382z4 = (Z382z4 & G482z4);
assign G482z4 = (~(Gzvvx4 & Gtnvx4));
assign Gtnvx4 = (~(N482z4 & U482z4));
assign U482z4 = (~(Tudvx4 & Jj9wx4));
assign N482z4 = (B582z4 & I582z4);
assign I582z4 = (~(Vb9wx4 & P582z4));
assign P582z4 = (~(W582z4 & D682z4));
assign D682z4 = (K682z4 & R682z4);
assign R682z4 = (Y682z4 & F782z4);
assign F782z4 = (~(vis_r14_o[24] & Zd9wx4));
assign Y682z4 = (M782z4 & T782z4);
assign T782z4 = (~(vis_psp_o[22] & Ue9wx4));
assign M782z4 = (~(vis_msp_o[22] & Bf9wx4));
assign K682z4 = (A882z4 & H882z4);
assign H882z4 = (~(vis_r12_o[24] & Wf9wx4));
assign A882z4 = (~(vis_r11_o[24] & Dg9wx4));
assign W582z4 = (O882z4 & V882z4);
assign V882z4 = (C982z4 & J982z4);
assign J982z4 = (~(vis_r10_o[24] & Mh9wx4));
assign C982z4 = (~(vis_r9_o[24] & Th9wx4));
assign O882z4 = (Mnvwx4 & Q982z4);
assign Q982z4 = (~(vis_r8_o[24] & Oi9wx4));
assign B582z4 = (~(Ewdvx4 & Qj9wx4));
assign Z382z4 = (~(Dmh2z4[24] & K1wvx4));
assign haddr_o[23] = (!Y92wx4);
assign Y92wx4 = (X982z4 & Ea82z4);
assign Ea82z4 = (~(Ykh2z4[22] & Mrsvx4));
assign X982z4 = (La82z4 & Sa82z4);
assign Sa82z4 = (~(Gzvvx4 & Ntnvx4));
assign Ntnvx4 = (~(Za82z4 & Gb82z4));
assign Gb82z4 = (~(Itdvx4 & Jj9wx4));
assign Za82z4 = (Nb82z4 & Ub82z4);
assign Ub82z4 = (~(Vb9wx4 & Bc82z4));
assign Bc82z4 = (~(Ic82z4 & Pc82z4));
assign Pc82z4 = (Wc82z4 & Dd82z4);
assign Dd82z4 = (Kd82z4 & Rd82z4);
assign Rd82z4 = (~(vis_r14_o[23] & Zd9wx4));
assign Kd82z4 = (Yd82z4 & Fe82z4);
assign Fe82z4 = (~(vis_psp_o[21] & Ue9wx4));
assign Yd82z4 = (~(vis_msp_o[21] & Bf9wx4));
assign Wc82z4 = (Me82z4 & Te82z4);
assign Te82z4 = (~(vis_r12_o[23] & Wf9wx4));
assign Me82z4 = (~(vis_r11_o[23] & Dg9wx4));
assign Ic82z4 = (Af82z4 & Hf82z4);
assign Hf82z4 = (Of82z4 & Vf82z4);
assign Vf82z4 = (~(vis_r10_o[23] & Mh9wx4));
assign Of82z4 = (~(vis_r9_o[23] & Th9wx4));
assign Af82z4 = (Icxwx4 & Cg82z4);
assign Cg82z4 = (~(vis_r8_o[23] & Oi9wx4));
assign Nb82z4 = (~(Tudvx4 & Qj9wx4));
assign La82z4 = (~(Dmh2z4[23] & K1wvx4));
assign haddr_o[22] = (!C70wx4);
assign C70wx4 = (Jg82z4 & Qg82z4);
assign Qg82z4 = (~(Ykh2z4[21] & Mrsvx4));
assign Jg82z4 = (Xg82z4 & Eh82z4);
assign Eh82z4 = (~(Gzvvx4 & Utnvx4));
assign Utnvx4 = (!N90wx4);
assign N90wx4 = (Lh82z4 & Sh82z4);
assign Sh82z4 = (~(Vb9wx4 & Zh82z4));
assign Zh82z4 = (~(Gi82z4 & Ni82z4));
assign Ni82z4 = (Ui82z4 & Bj82z4);
assign Bj82z4 = (Ij82z4 & Pj82z4);
assign Pj82z4 = (~(Zd9wx4 & vis_r14_o[22]));
assign Ij82z4 = (Wj82z4 & Dk82z4);
assign Dk82z4 = (~(Ue9wx4 & vis_psp_o[20]));
assign Wj82z4 = (~(Bf9wx4 & vis_msp_o[20]));
assign Ui82z4 = (Kk82z4 & Rk82z4);
assign Rk82z4 = (~(Wf9wx4 & vis_r12_o[22]));
assign Kk82z4 = (~(Dg9wx4 & vis_r11_o[22]));
assign Gi82z4 = (Yk82z4 & Fl82z4);
assign Fl82z4 = (Ml82z4 & Tl82z4);
assign Tl82z4 = (~(Mh9wx4 & vis_r10_o[22]));
assign Ml82z4 = (~(Th9wx4 & vis_r9_o[22]));
assign Yk82z4 = (G4qwx4 & Am82z4);
assign Am82z4 = (~(Oi9wx4 & vis_r8_o[22]));
assign Lh82z4 = (Hm82z4 & Om82z4);
assign Om82z4 = (~(Xrdvx4 & Jj9wx4));
assign Hm82z4 = (~(Qj9wx4 & Itdvx4));
assign Xg82z4 = (~(Dmh2z4[22] & K1wvx4));
assign haddr_o[21] = (!Fc0wx4);
assign Fc0wx4 = (Vm82z4 & Cn82z4);
assign Cn82z4 = (~(Ykh2z4[20] & Mrsvx4));
assign Vm82z4 = (Jn82z4 & Qn82z4);
assign Qn82z4 = (~(Gzvvx4 & Bunvx4));
assign Bunvx4 = (!Lf0wx4);
assign Lf0wx4 = (Xn82z4 & Eo82z4);
assign Eo82z4 = (~(Vb9wx4 & Lo82z4));
assign Lo82z4 = (~(So82z4 & Zo82z4));
assign Zo82z4 = (Gp82z4 & Np82z4);
assign Np82z4 = (Up82z4 & Bq82z4);
assign Bq82z4 = (~(Zd9wx4 & vis_r14_o[21]));
assign Up82z4 = (Iq82z4 & Pq82z4);
assign Pq82z4 = (~(Ue9wx4 & vis_psp_o[19]));
assign Iq82z4 = (~(Bf9wx4 & vis_msp_o[19]));
assign Gp82z4 = (Wq82z4 & Dr82z4);
assign Dr82z4 = (~(Wf9wx4 & vis_r12_o[21]));
assign Wq82z4 = (~(Dg9wx4 & vis_r11_o[21]));
assign So82z4 = (Kr82z4 & Rr82z4);
assign Rr82z4 = (Yr82z4 & Fs82z4);
assign Fs82z4 = (~(Mh9wx4 & vis_r10_o[21]));
assign Yr82z4 = (~(Th9wx4 & vis_r9_o[21]));
assign Kr82z4 = (D9uwx4 & Ms82z4);
assign Ms82z4 = (~(Oi9wx4 & vis_r8_o[21]));
assign Xn82z4 = (Ts82z4 & At82z4);
assign At82z4 = (~(Mqdvx4 & Jj9wx4));
assign Ts82z4 = (~(Qj9wx4 & Xrdvx4));
assign Jn82z4 = (~(Dmh2z4[21] & K1wvx4));
assign haddr_o[20] = (!Ug0wx4);
assign Ug0wx4 = (Ht82z4 & Ot82z4);
assign Ot82z4 = (~(Ykh2z4[19] & Mrsvx4));
assign Ht82z4 = (Vt82z4 & Cu82z4);
assign Cu82z4 = (~(Gzvvx4 & Iunvx4));
assign Iunvx4 = (!Fj0wx4);
assign Fj0wx4 = (Ju82z4 & Qu82z4);
assign Qu82z4 = (~(Vb9wx4 & Xu82z4));
assign Xu82z4 = (~(Ev82z4 & Lv82z4));
assign Lv82z4 = (Sv82z4 & Zv82z4);
assign Zv82z4 = (Gw82z4 & Nw82z4);
assign Nw82z4 = (~(Zd9wx4 & vis_r14_o[20]));
assign Gw82z4 = (Uw82z4 & Bx82z4);
assign Bx82z4 = (~(Ue9wx4 & vis_psp_o[18]));
assign Uw82z4 = (~(Bf9wx4 & vis_msp_o[18]));
assign Sv82z4 = (Ix82z4 & Px82z4);
assign Px82z4 = (~(Wf9wx4 & vis_r12_o[20]));
assign Ix82z4 = (~(Dg9wx4 & vis_r11_o[20]));
assign Ev82z4 = (Wx82z4 & Dy82z4);
assign Dy82z4 = (Ky82z4 & Ry82z4);
assign Ry82z4 = (~(Mh9wx4 & vis_r10_o[20]));
assign Ky82z4 = (~(Th9wx4 & vis_r9_o[20]));
assign Wx82z4 = (Dmvwx4 & Yy82z4);
assign Yy82z4 = (~(Oi9wx4 & vis_r8_o[20]));
assign Ju82z4 = (Fz82z4 & Mz82z4);
assign Mz82z4 = (~(Bpdvx4 & Jj9wx4));
assign Fz82z4 = (~(Qj9wx4 & Mqdvx4));
assign Vt82z4 = (~(Dmh2z4[20] & K1wvx4));
assign haddr_o[1] = (~(Y162z4 | Loyvx4));
assign Loyvx4 = (!T50wx4);
assign T50wx4 = (~(Tz82z4 & A092z4));
assign A092z4 = (~(Dmh2z4[1] & K1wvx4));
assign Tz82z4 = (H092z4 & O092z4);
assign O092z4 = (~(Mrsvx4 & V092z4));
assign V092z4 = (~(vis_pc_o[0] ^ Zorvx4));
assign H092z4 = (~(Gzvvx4 & Punvx4));
assign Punvx4 = (~(C192z4 & J192z4));
assign J192z4 = (~(Kycvx4 & Jj9wx4));
assign C192z4 = (Q192z4 & X192z4);
assign X192z4 = (~(Vb9wx4 & E292z4));
assign E292z4 = (~(L292z4 & S292z4));
assign S292z4 = (Z292z4 & G392z4);
assign G392z4 = (N392z4 & U392z4);
assign U392z4 = (~(vis_r14_o[1] & Zd9wx4));
assign N392z4 = (~(vis_r12_o[1] & Wf9wx4));
assign Z292z4 = (B492z4 & I492z4);
assign I492z4 = (~(vis_r11_o[1] & Dg9wx4));
assign B492z4 = (~(vis_r10_o[1] & Mh9wx4));
assign L292z4 = (P492z4 & Duuwx4);
assign P492z4 = (W492z4 & D592z4);
assign D592z4 = (~(vis_r9_o[1] & Th9wx4));
assign W492z4 = (~(vis_r8_o[1] & Oi9wx4));
assign Q192z4 = (~(Uzcvx4 & Qj9wx4));
assign haddr_o[19] = (!Ql0wx4);
assign Ql0wx4 = (K592z4 & R592z4);
assign R592z4 = (~(Ykh2z4[18] & Mrsvx4));
assign K592z4 = (Y592z4 & F692z4);
assign F692z4 = (~(Gzvvx4 & Wunvx4));
assign Wunvx4 = (!Wo0wx4);
assign Wo0wx4 = (M692z4 & T692z4);
assign T692z4 = (~(Vb9wx4 & A792z4));
assign A792z4 = (~(H792z4 & O792z4));
assign O792z4 = (V792z4 & C892z4);
assign C892z4 = (J892z4 & Q892z4);
assign Q892z4 = (~(Zd9wx4 & vis_r14_o[19]));
assign J892z4 = (X892z4 & E992z4);
assign E992z4 = (~(Ue9wx4 & vis_psp_o[17]));
assign X892z4 = (~(Bf9wx4 & vis_msp_o[17]));
assign V792z4 = (L992z4 & S992z4);
assign S992z4 = (~(Wf9wx4 & vis_r12_o[19]));
assign L992z4 = (~(Dg9wx4 & vis_r11_o[19]));
assign H792z4 = (Z992z4 & Ga92z4);
assign Ga92z4 = (Na92z4 & Ua92z4);
assign Ua92z4 = (~(Mh9wx4 & vis_r10_o[19]));
assign Na92z4 = (~(Th9wx4 & vis_r9_o[19]));
assign Z992z4 = (Bjxwx4 & Bb92z4);
assign Bb92z4 = (~(Oi9wx4 & vis_r8_o[19]));
assign M692z4 = (Ib92z4 & Pb92z4);
assign Pb92z4 = (~(Qndvx4 & Jj9wx4));
assign Ib92z4 = (~(Qj9wx4 & Bpdvx4));
assign Y592z4 = (~(Dmh2z4[19] & K1wvx4));
assign haddr_o[18] = (!Fq0wx4);
assign Fq0wx4 = (Wb92z4 & Dc92z4);
assign Dc92z4 = (~(Ykh2z4[17] & Mrsvx4));
assign Wb92z4 = (Kc92z4 & Rc92z4);
assign Rc92z4 = (~(Gzvvx4 & Dvnvx4));
assign Dvnvx4 = (!Qs0wx4);
assign Qs0wx4 = (Yc92z4 & Fd92z4);
assign Fd92z4 = (~(Vb9wx4 & Md92z4));
assign Md92z4 = (~(Td92z4 & Ae92z4));
assign Ae92z4 = (He92z4 & Oe92z4);
assign Oe92z4 = (Ve92z4 & Cf92z4);
assign Cf92z4 = (~(Zd9wx4 & vis_r14_o[18]));
assign Ve92z4 = (Jf92z4 & Qf92z4);
assign Qf92z4 = (~(Ue9wx4 & vis_psp_o[16]));
assign Jf92z4 = (~(Bf9wx4 & vis_msp_o[16]));
assign He92z4 = (Xf92z4 & Eg92z4);
assign Eg92z4 = (~(Wf9wx4 & vis_r12_o[18]));
assign Xf92z4 = (~(Dg9wx4 & vis_r11_o[18]));
assign Td92z4 = (Lg92z4 & Sg92z4);
assign Sg92z4 = (Zg92z4 & Gh92z4);
assign Gh92z4 = (~(Mh9wx4 & vis_r10_o[18]));
assign Zg92z4 = (~(Th9wx4 & vis_r9_o[18]));
assign Lg92z4 = (H1qwx4 & Nh92z4);
assign Nh92z4 = (~(Oi9wx4 & vis_r8_o[18]));
assign Yc92z4 = (Uh92z4 & Bi92z4);
assign Bi92z4 = (~(Fmdvx4 & Jj9wx4));
assign Uh92z4 = (~(Qj9wx4 & Qndvx4));
assign Kc92z4 = (~(Dmh2z4[18] & K1wvx4));
assign haddr_o[17] = (!Bv0wx4);
assign Bv0wx4 = (Ii92z4 & Pi92z4);
assign Pi92z4 = (~(Ykh2z4[16] & Mrsvx4));
assign Ii92z4 = (Wi92z4 & Dj92z4);
assign Dj92z4 = (~(Gzvvx4 & Kvnvx4));
assign Kvnvx4 = (!Hy0wx4);
assign Hy0wx4 = (Kj92z4 & Rj92z4);
assign Rj92z4 = (~(Vb9wx4 & Yj92z4));
assign Yj92z4 = (~(Fk92z4 & Mk92z4));
assign Mk92z4 = (Tk92z4 & Al92z4);
assign Al92z4 = (Hl92z4 & Ol92z4);
assign Ol92z4 = (~(Zd9wx4 & vis_r14_o[17]));
assign Hl92z4 = (Vl92z4 & Cm92z4);
assign Cm92z4 = (~(Ue9wx4 & vis_psp_o[15]));
assign Vl92z4 = (~(Bf9wx4 & vis_msp_o[15]));
assign Tk92z4 = (Jm92z4 & Qm92z4);
assign Qm92z4 = (~(Wf9wx4 & vis_r12_o[17]));
assign Jm92z4 = (~(Dg9wx4 & vis_r11_o[17]));
assign Fk92z4 = (Xm92z4 & En92z4);
assign En92z4 = (Ln92z4 & Sn92z4);
assign Sn92z4 = (~(Mh9wx4 & vis_r10_o[17]));
assign Ln92z4 = (~(Th9wx4 & vis_r9_o[17]));
assign Xm92z4 = (Xcuwx4 & Zn92z4);
assign Zn92z4 = (~(Oi9wx4 & vis_r8_o[17]));
assign Kj92z4 = (Go92z4 & No92z4);
assign No92z4 = (~(Ukdvx4 & Jj9wx4));
assign Go92z4 = (~(Qj9wx4 & Fmdvx4));
assign Wi92z4 = (~(Dmh2z4[17] & K1wvx4));
assign haddr_o[16] = (!Vpovx4);
assign Vpovx4 = (Uo92z4 & Bp92z4);
assign Bp92z4 = (~(Ykh2z4[15] & Mrsvx4));
assign Uo92z4 = (Ip92z4 & Pp92z4);
assign Pp92z4 = (~(Gzvvx4 & Rvnvx4));
assign Rvnvx4 = (!U11wx4);
assign U11wx4 = (Wp92z4 & Dq92z4);
assign Dq92z4 = (~(Vb9wx4 & Kq92z4));
assign Kq92z4 = (~(Rq92z4 & Yq92z4));
assign Yq92z4 = (Fr92z4 & Mr92z4);
assign Mr92z4 = (Tr92z4 & As92z4);
assign As92z4 = (~(Zd9wx4 & vis_r14_o[16]));
assign Tr92z4 = (Hs92z4 & Os92z4);
assign Os92z4 = (~(Ue9wx4 & vis_psp_o[14]));
assign Hs92z4 = (~(Bf9wx4 & vis_msp_o[14]));
assign Fr92z4 = (Vs92z4 & Ct92z4);
assign Ct92z4 = (~(Wf9wx4 & vis_r12_o[16]));
assign Vs92z4 = (~(Dg9wx4 & vis_r11_o[16]));
assign Rq92z4 = (Jt92z4 & Qt92z4);
assign Qt92z4 = (Xt92z4 & Eu92z4);
assign Eu92z4 = (~(Mh9wx4 & vis_r10_o[16]));
assign Xt92z4 = (~(Th9wx4 & vis_r9_o[16]));
assign Jt92z4 = (Nrvwx4 & Lu92z4);
assign Lu92z4 = (~(Oi9wx4 & vis_r8_o[16]));
assign Wp92z4 = (Su92z4 & Zu92z4);
assign Zu92z4 = (~(Jjdvx4 & Jj9wx4));
assign Su92z4 = (~(Qj9wx4 & Ukdvx4));
assign Ip92z4 = (~(Dmh2z4[16] & K1wvx4));
assign haddr_o[14] = (~(Gv92z4 & Nv92z4));
assign Nv92z4 = (~(Ykh2z4[13] & Mrsvx4));
assign Gv92z4 = (Uv92z4 & Bw92z4);
assign Bw92z4 = (~(Gzvvx4 & Fwnvx4));
assign Fwnvx4 = (!C61wx4);
assign C61wx4 = (Iw92z4 & Pw92z4);
assign Pw92z4 = (~(Vb9wx4 & Ww92z4));
assign Ww92z4 = (~(Dx92z4 & Kx92z4));
assign Kx92z4 = (Rx92z4 & Yx92z4);
assign Yx92z4 = (Fy92z4 & My92z4);
assign My92z4 = (~(Zd9wx4 & vis_r14_o[14]));
assign Fy92z4 = (Ty92z4 & Az92z4);
assign Az92z4 = (~(Ue9wx4 & vis_psp_o[12]));
assign Ty92z4 = (~(Bf9wx4 & vis_msp_o[12]));
assign Rx92z4 = (Hz92z4 & Oz92z4);
assign Oz92z4 = (~(Wf9wx4 & vis_r12_o[14]));
assign Hz92z4 = (~(Dg9wx4 & vis_r11_o[14]));
assign Dx92z4 = (Vz92z4 & C0a2z4);
assign C0a2z4 = (J0a2z4 & Q0a2z4);
assign Q0a2z4 = (~(Mh9wx4 & vis_r10_o[14]));
assign J0a2z4 = (~(Th9wx4 & vis_r9_o[14]));
assign Vz92z4 = (Hmqwx4 & X0a2z4);
assign X0a2z4 = (~(Oi9wx4 & vis_r8_o[14]));
assign Iw92z4 = (E1a2z4 & L1a2z4);
assign L1a2z4 = (~(Ngdvx4 & Jj9wx4));
assign E1a2z4 = (~(Qj9wx4 & Yhdvx4));
assign Uv92z4 = (~(Dmh2z4[14] & K1wvx4));
assign haddr_o[13] = (~(S1a2z4 & Z1a2z4));
assign Z1a2z4 = (~(Ykh2z4[12] & Mrsvx4));
assign S1a2z4 = (G2a2z4 & N2a2z4);
assign N2a2z4 = (~(Gzvvx4 & Mwnvx4));
assign Mwnvx4 = (!Ra1wx4);
assign Ra1wx4 = (U2a2z4 & B3a2z4);
assign B3a2z4 = (~(Vb9wx4 & I3a2z4));
assign I3a2z4 = (~(P3a2z4 & W3a2z4));
assign W3a2z4 = (D4a2z4 & K4a2z4);
assign K4a2z4 = (R4a2z4 & Y4a2z4);
assign Y4a2z4 = (~(Zd9wx4 & vis_r14_o[13]));
assign R4a2z4 = (F5a2z4 & M5a2z4);
assign M5a2z4 = (~(Ue9wx4 & vis_psp_o[11]));
assign F5a2z4 = (~(Bf9wx4 & vis_msp_o[11]));
assign D4a2z4 = (T5a2z4 & A6a2z4);
assign A6a2z4 = (~(Wf9wx4 & vis_r12_o[13]));
assign T5a2z4 = (~(Dg9wx4 & vis_r11_o[13]));
assign P3a2z4 = (H6a2z4 & O6a2z4);
assign O6a2z4 = (V6a2z4 & C7a2z4);
assign C7a2z4 = (~(Mh9wx4 & vis_r10_o[13]));
assign V6a2z4 = (~(Th9wx4 & vis_r9_o[13]));
assign H6a2z4 = (Zkuwx4 & J7a2z4);
assign J7a2z4 = (~(Oi9wx4 & vis_r8_o[13]));
assign U2a2z4 = (Q7a2z4 & X7a2z4);
assign X7a2z4 = (~(Cfdvx4 & Jj9wx4));
assign Q7a2z4 = (~(Qj9wx4 & Ngdvx4));
assign G2a2z4 = (~(Dmh2z4[13] & K1wvx4));
assign haddr_o[12] = (!Cqovx4);
assign Cqovx4 = (E8a2z4 & L8a2z4);
assign L8a2z4 = (~(Ykh2z4[11] & Mrsvx4));
assign E8a2z4 = (S8a2z4 & Z8a2z4);
assign Z8a2z4 = (~(Gzvvx4 & Twnvx4));
assign Twnvx4 = (!Pg1wx4);
assign Pg1wx4 = (G9a2z4 & N9a2z4);
assign N9a2z4 = (~(Vb9wx4 & U9a2z4));
assign U9a2z4 = (~(Baa2z4 & Iaa2z4));
assign Iaa2z4 = (Paa2z4 & Waa2z4);
assign Waa2z4 = (Dba2z4 & Kba2z4);
assign Kba2z4 = (~(Zd9wx4 & vis_r14_o[12]));
assign Dba2z4 = (Rba2z4 & Yba2z4);
assign Yba2z4 = (~(Ue9wx4 & vis_psp_o[10]));
assign Rba2z4 = (~(Bf9wx4 & vis_msp_o[10]));
assign Paa2z4 = (Fca2z4 & Mca2z4);
assign Mca2z4 = (~(Wf9wx4 & vis_r12_o[12]));
assign Fca2z4 = (~(Dg9wx4 & vis_r11_o[12]));
assign Baa2z4 = (Tca2z4 & Ada2z4);
assign Ada2z4 = (Hda2z4 & Oda2z4);
assign Oda2z4 = (~(Mh9wx4 & vis_r10_o[12]));
assign Hda2z4 = (~(Th9wx4 & vis_r9_o[12]));
assign Tca2z4 = (H2wwx4 & Vda2z4);
assign Vda2z4 = (~(Oi9wx4 & vis_r8_o[12]));
assign G9a2z4 = (Cea2z4 & Jea2z4);
assign Jea2z4 = (~(Rddvx4 & Jj9wx4));
assign Cea2z4 = (~(Qj9wx4 & Cfdvx4));
assign S8a2z4 = (~(Dmh2z4[12] & K1wvx4));
assign haddr_o[10] = (!Jxovx4);
assign Jxovx4 = (Qea2z4 & Xea2z4);
assign Xea2z4 = (~(Ykh2z4[9] & Mrsvx4));
assign Qea2z4 = (Efa2z4 & Lfa2z4);
assign Lfa2z4 = (~(Gzvvx4 & Hxnvx4));
assign Hxnvx4 = (~(Sfa2z4 & Zfa2z4));
assign Zfa2z4 = (~(Wadvx4 & Jj9wx4));
assign Sfa2z4 = (Gga2z4 & Nga2z4);
assign Nga2z4 = (~(Vb9wx4 & Uga2z4));
assign Uga2z4 = (~(Bha2z4 & Iha2z4));
assign Iha2z4 = (Pha2z4 & Wha2z4);
assign Wha2z4 = (Dia2z4 & Kia2z4);
assign Kia2z4 = (~(vis_r14_o[10] & Zd9wx4));
assign Dia2z4 = (Ria2z4 & Yia2z4);
assign Yia2z4 = (~(vis_psp_o[8] & Ue9wx4));
assign Ue9wx4 = (Fja2z4 & Mja2z4);
assign Fja2z4 = (~(Tja2z4 | Ta2wx4));
assign Ta2wx4 = (!O7evx4);
assign Ria2z4 = (~(vis_msp_o[8] & Bf9wx4));
assign Bf9wx4 = (Aka2z4 & Mja2z4);
assign Aka2z4 = (~(Tja2z4 | O7evx4));
assign Pha2z4 = (Hka2z4 & Oka2z4);
assign Oka2z4 = (~(vis_r12_o[10] & Wf9wx4));
assign Hka2z4 = (~(vis_r11_o[10] & Dg9wx4));
assign Bha2z4 = (Vka2z4 & Cla2z4);
assign Cla2z4 = (Jla2z4 & Qla2z4);
assign Qla2z4 = (~(vis_r10_o[10] & Mh9wx4));
assign Jla2z4 = (~(vis_r9_o[10] & Th9wx4));
assign Vka2z4 = (Pjqwx4 & Xla2z4);
assign Xla2z4 = (~(vis_r8_o[10] & Oi9wx4));
assign Gga2z4 = (~(Gcdvx4 & Qj9wx4));
assign Efa2z4 = (~(Dmh2z4[10] & K1wvx4));
assign haddr_o[0] = (~(Ema2z4 | Y162z4));
assign Y162z4 = (~(Qr42z4 & It52z4));
assign It52z4 = (~(Lma2z4 & Sma2z4));
assign Sma2z4 = (Wpsvx4 & Z5pvx4);
assign Z5pvx4 = (Zma2z4 & Gna2z4);
assign Gna2z4 = (~(Rkgvx4 & Nna2z4));
assign Nna2z4 = (~(Ik4wx4 & Una2z4));
assign Ik4wx4 = (Boa2z4 & Ioa2z4);
assign Ioa2z4 = (Poa2z4 & Woa2z4);
assign Woa2z4 = (~(Dpa2z4 & Kpa2z4));
assign Kpa2z4 = (~(J43wx4 | C34wx4));
assign C34wx4 = (Rpa2z4 & Ypa2z4);
assign Ypa2z4 = (~(Fqa2z4 & Xtywx4));
assign Xtywx4 = (~(Mqa2z4 & Tqa2z4));
assign Tqa2z4 = (Ara2z4 & Hra2z4);
assign Hra2z4 = (Ora2z4 & Vra2z4);
assign Vra2z4 = (Csa2z4 & Kvuvx4);
assign Csa2z4 = (~(Jsa2z4 | Qsa2z4));
assign Qsa2z4 = (!Yauvx4);
assign Ora2z4 = (~(K9ovx4 | Jruvx4));
assign Ara2z4 = (Xsa2z4 & Eta2z4);
assign Eta2z4 = (Lta2z4 & Ruvvx4);
assign Lta2z4 = (~(Sta2z4 | Zta2z4));
assign Xsa2z4 = (~(Pguvx4 | Gua2z4));
assign Gua2z4 = (!Ckuvx4);
assign Mqa2z4 = (Nua2z4 & Uua2z4);
assign Uua2z4 = (Bva2z4 & Iva2z4);
assign Iva2z4 = (Pva2z4 & Mhvvx4);
assign Pva2z4 = (~(Wva2z4 | Dwa2z4));
assign Dwa2z4 = (!K9vvx4);
assign Bva2z4 = (~(Oxuvx4 | Kwa2z4));
assign Nua2z4 = (Rwa2z4 & Ywa2z4);
assign Ywa2z4 = (~(Fxa2z4 | Mxa2z4));
assign Rwa2z4 = (~(Douvx4 | Txa2z4));
assign Fqa2z4 = (~(Aya2z4 & Hya2z4));
assign Hya2z4 = (~(Uth2z4[1] & Oya2z4));
assign Oya2z4 = (~(Vya2z4 & Vsywx4));
assign Aya2z4 = (Vsywx4 | Vya2z4);
assign Vya2z4 = (Iwywx4 & Luywx4);
assign Luywx4 = (~(Cza2z4 & Jza2z4));
assign Jza2z4 = (Qza2z4 & Xza2z4);
assign Xza2z4 = (E0b2z4 & L0b2z4);
assign L0b2z4 = (S0b2z4 & Z0b2z4);
assign Z0b2z4 = (~(Zuh2z4[8] & Oxuvx4));
assign S0b2z4 = (G1b2z4 & N1b2z4);
assign N1b2z4 = (Vgpwx4 | Hpvvx4);
assign Vgpwx4 = (!Txh2z4[0]);
assign G1b2z4 = (J3pwx4 | Uevvx4);
assign J3pwx4 = (!Zuh2z4[18]);
assign E0b2z4 = (U1b2z4 & B2b2z4);
assign B2b2z4 = (~(Zuh2z4[24] & Kwa2z4));
assign U1b2z4 = (Tmpwx4 | Mhvvx4);
assign Tmpwx4 = (!Zuh2z4[16]);
assign Qza2z4 = (I2b2z4 & P2b2z4);
assign P2b2z4 = (W2b2z4 & D3b2z4);
assign D3b2z4 = (Chpwx4 | K9vvx4);
assign Chpwx4 = (!Zuh2z4[22]);
assign W2b2z4 = (K3b2z4 & R3b2z4);
assign R3b2z4 = (Zxowx4 | Ccvvx4);
assign Zxowx4 = (!Zuh2z4[20]);
assign K3b2z4 = (Sipwx4 | Fpuvx4);
assign Sipwx4 = (!Zuh2z4[14]);
assign I2b2z4 = (Y3b2z4 & F4b2z4);
assign F4b2z4 = (Njpwx4 | Khuvx4);
assign Njpwx4 = (!Zuh2z4[6]);
assign Y3b2z4 = (Uyowx4 | Ckuvx4);
assign Uyowx4 = (!Zuh2z4[4]);
assign Cza2z4 = (M4b2z4 & T4b2z4);
assign T4b2z4 = (A5b2z4 & H5b2z4);
assign H5b2z4 = (O5b2z4 & V5b2z4);
assign V5b2z4 = (Sxowx4 | Rnvvx4);
assign Sxowx4 = (!Psh2z4[0]);
assign O5b2z4 = (C6b2z4 & J6b2z4);
assign J6b2z4 = (O9pwx4 | Ruvvx4);
assign O9pwx4 = (!Zuh2z4[2]);
assign C6b2z4 = (Iwywx4 | Oivvx4);
assign Oivvx4 = (!Sta2z4);
assign A5b2z4 = (Q6b2z4 & X6b2z4);
assign X6b2z4 = (Onpwx4 | Taovx4);
assign Onpwx4 = (!Zuh2z4[0]);
assign Q6b2z4 = (~(Zuh2z4[12] & Jruvx4));
assign M4b2z4 = (E7b2z4 & L7b2z4);
assign L7b2z4 = (S7b2z4 & Z7b2z4);
assign Z7b2z4 = (R7pwx4 | Kvuvx4);
assign R7pwx4 = (!Zuh2z4[10]);
assign S7b2z4 = (Lipwx4 | G8uvx4);
assign Lipwx4 = (!Zuh2z4[30]);
assign E7b2z4 = (G8b2z4 & N8b2z4);
assign N8b2z4 = (Xwowx4 | Jxvvx4);
assign Xwowx4 = (!Zuh2z4[28]);
assign G8b2z4 = (D7pwx4 | Yauvx4);
assign D7pwx4 = (!Zuh2z4[26]);
assign Iwywx4 = (!Uth2z4[0]);
assign Vsywx4 = (~(U8b2z4 & B9b2z4));
assign B9b2z4 = (I9b2z4 & P9b2z4);
assign P9b2z4 = (W9b2z4 & Dab2z4);
assign Dab2z4 = (Kab2z4 & Rab2z4);
assign Rab2z4 = (Wbywx4 | Hpvvx4);
assign Hpvvx4 = (!Fxa2z4);
assign Fxa2z4 = (Yab2z4 & Fbb2z4);
assign Wbywx4 = (!Txh2z4[1]);
assign Kab2z4 = (Mbb2z4 & Tbb2z4);
assign Tbb2z4 = (Iqxwx4 | Ruvvx4);
assign Ruvvx4 = (~(Acb2z4 & Hcb2z4));
assign Acb2z4 = (Ocb2z4 & T0rvx4);
assign Iqxwx4 = (!Zuh2z4[3]);
assign Mbb2z4 = (J9xwx4 | Ccvvx4);
assign Ccvvx4 = (!Wva2z4);
assign Wva2z4 = (Vcb2z4 & Cdb2z4);
assign J9xwx4 = (!Zuh2z4[21]);
assign W9b2z4 = (Jdb2z4 & Qdb2z4);
assign Qdb2z4 = (Xnxwx4 | Kvuvx4);
assign Kvuvx4 = (!Iuuvx4);
assign Iuuvx4 = (Ocb2z4 & Xdb2z4);
assign Xnxwx4 = (!Zuh2z4[11]);
assign Jdb2z4 = (~(Uth2z4[1] & Sta2z4));
assign Sta2z4 = (Eeb2z4 & Fbb2z4);
assign I9b2z4 = (Leb2z4 & Seb2z4);
assign Seb2z4 = (Zeb2z4 & Gfb2z4);
assign Gfb2z4 = (Eaxwx4 | Esuvx4);
assign Esuvx4 = (!Jruvx4);
assign Jruvx4 = (Nfb2z4 & Ocb2z4);
assign Eaxwx4 = (!Zuh2z4[13]);
assign Zeb2z4 = (Ufb2z4 & Bgb2z4);
assign Bgb2z4 = (C9xwx4 | Rnvvx4);
assign Rnvvx4 = (!Zta2z4);
assign Zta2z4 = (Nfb2z4 & Fbb2z4);
assign Fbb2z4 = (Igb2z4 & vis_ipsr_o[3]);
assign Nfb2z4 = (Pgb2z4 & Gxqvx4);
assign C9xwx4 = (!Psh2z4[1]);
assign Ufb2z4 = (C2xwx4 | Taovx4);
assign Taovx4 = (!K9ovx4);
assign K9ovx4 = (Wgb2z4 & Ocb2z4);
assign C2xwx4 = (!Zuh2z4[1]);
assign Leb2z4 = (Dhb2z4 & Khb2z4);
assign Khb2z4 = (Fdywx4 | K9vvx4);
assign K9vvx4 = (~(Eeb2z4 & Cdb2z4));
assign Fdywx4 = (!Zuh2z4[23]);
assign Dhb2z4 = (Jfywx4 | Fpuvx4);
assign Fpuvx4 = (!Douvx4);
assign Douvx4 = (Yab2z4 & Ocb2z4);
assign Yab2z4 = (Pgb2z4 & vis_ipsr_o[0]);
assign Jfywx4 = (!Zuh2z4[15]);
assign U8b2z4 = (Rhb2z4 & Yhb2z4);
assign Yhb2z4 = (Fib2z4 & Mib2z4);
assign Mib2z4 = (Tib2z4 & Ajb2z4);
assign Ajb2z4 = (A1xwx4 | Ulvvx4);
assign Ulvvx4 = (!Kwa2z4);
assign Kwa2z4 = (Hjb2z4 & Cdb2z4);
assign A1xwx4 = (!Zuh2z4[25]);
assign Tib2z4 = (Ojb2z4 & Vjb2z4);
assign Vjb2z4 = (V1xwx4 | Qyuvx4);
assign Qyuvx4 = (!Oxuvx4);
assign Oxuvx4 = (Hjb2z4 & Ocb2z4);
assign Hjb2z4 = (vis_ipsr_o[2] & Ckb2z4);
assign V1xwx4 = (!Zuh2z4[9]);
assign Ojb2z4 = (Omxwx4 | Uevvx4);
assign Uevvx4 = (!Mxa2z4);
assign Mxa2z4 = (Jkb2z4 & Hcb2z4);
assign Jkb2z4 = (Cdb2z4 & T0rvx4);
assign Omxwx4 = (!Zuh2z4[19]);
assign Fib2z4 = (Qkb2z4 & Xkb2z4);
assign Xkb2z4 = (T0xwx4 | Mhvvx4);
assign Mhvvx4 = (~(Wgb2z4 & Cdb2z4));
assign T0xwx4 = (!Zuh2z4[17]);
assign Qkb2z4 = (Xfywx4 | Khuvx4);
assign Khuvx4 = (!Pguvx4);
assign Pguvx4 = (Eeb2z4 & Ocb2z4);
assign Eeb2z4 = (Hcb2z4 & vis_ipsr_o[1]);
assign Hcb2z4 = (vis_ipsr_o[0] & Xkuvx4);
assign Xfywx4 = (!Zuh2z4[7]);
assign Rhb2z4 = (Elb2z4 & Llb2z4);
assign Llb2z4 = (Slb2z4 & Zlb2z4);
assign Zlb2z4 = (Laxwx4 | Ckuvx4);
assign Ckuvx4 = (~(Vcb2z4 & Ocb2z4));
assign Ocb2z4 = (Gmb2z4 & vis_ipsr_o[4]);
assign Gmb2z4 = (~(vis_ipsr_o[3] | vis_ipsr_o[5]));
assign Vcb2z4 = (Nmb2z4 & vis_ipsr_o[1]);
assign Nmb2z4 = (~(vis_ipsr_o[0] | vis_ipsr_o[2]));
assign Laxwx4 = (!Zuh2z4[5]);
assign Slb2z4 = (H8xwx4 | Jxvvx4);
assign Jxvvx4 = (!Txa2z4);
assign Txa2z4 = (Umb2z4 & Pgb2z4);
assign Umb2z4 = (Cdb2z4 & Gxqvx4);
assign H8xwx4 = (!Zuh2z4[29]);
assign Elb2z4 = (Bnb2z4 & Inb2z4);
assign Inb2z4 = (Tlxwx4 | Yauvx4);
assign Yauvx4 = (~(Xdb2z4 & Cdb2z4));
assign Xdb2z4 = (Pnb2z4 & vis_ipsr_o[2]);
assign Pnb2z4 = (~(Gxqvx4 | vis_ipsr_o[1]));
assign Tlxwx4 = (!Zuh2z4[27]);
assign Bnb2z4 = (Tdywx4 | G8uvx4);
assign G8uvx4 = (!Jsa2z4);
assign Jsa2z4 = (Wnb2z4 & Pgb2z4);
assign Pgb2z4 = (vis_ipsr_o[2] & vis_ipsr_o[1]);
assign Wnb2z4 = (Cdb2z4 & vis_ipsr_o[0]);
assign Cdb2z4 = (Dob2z4 & vis_ipsr_o[4]);
assign Dob2z4 = (~(Lzuvx4 | vis_ipsr_o[5]));
assign Tdywx4 = (!Zuh2z4[31]);
assign Rpa2z4 = (~(Ye4wx4 | vis_primask_o));
assign Ye4wx4 = (Kob2z4 & Rob2z4);
assign Kob2z4 = (~(T0rvx4 | vis_ipsr_o[2]));
assign Dpa2z4 = (E44wx4 & Z7fwx4);
assign Poa2z4 = (~(Yob2z4 & D8hwx4));
assign D8hwx4 = (Fpb2z4 & C2yvx4);
assign Fpb2z4 = (~(Tv2wx4 | Fpfwx4));
assign Yob2z4 = (Pcyvx4 & Mpb2z4);
assign Mpb2z4 = (!W7hwx4);
assign Boa2z4 = (Wpsvx4 & Tpb2z4);
assign Tpb2z4 = (~(Bk4wx4 & Aqb2z4));
assign Aqb2z4 = (Hqb2z4 | Oqb2z4);
assign Oqb2z4 = (Xmsvx4 ? Lcpvx4 : Vqb2z4);
assign Lcpvx4 = (!Aj9vx4);
assign Vqb2z4 = (~(Ho8vx4 | Cf9vx4));
assign Hqb2z4 = (Mgwvx4 | O1jwx4);
assign Bk4wx4 = (Crb2z4 & Jrb2z4);
assign Jrb2z4 = (~(S4xvx4 | T93wx4));
assign Crb2z4 = (~(Fscwx4 | U4yvx4));
assign U4yvx4 = (!Rngwx4);
assign Zma2z4 = (Qrb2z4 & Xrb2z4);
assign Xrb2z4 = (~(Esb2z4 & Pcyvx4));
assign Esb2z4 = (Lsb2z4 & F3ovx4);
assign Lsb2z4 = (~(Ssb2z4 & Zsb2z4));
assign Zsb2z4 = (~(Gtb2z4 & Ntb2z4));
assign Ntb2z4 = (C2yvx4 & Rkgvx4);
assign Gtb2z4 = (~(Fscwx4 | Oedwx4));
assign Fscwx4 = (!D83wx4);
assign D83wx4 = (~(W5yvx4 | Dbgvx4));
assign Ssb2z4 = (~(Fqlwx4 & Nv6wx4));
assign Qrb2z4 = (~(Utb2z4 & P5yvx4));
assign Utb2z4 = (~(R7qvx4 | T93wx4));
assign Lma2z4 = (Bub2z4 & Ppsvx4);
assign Ppsvx4 = (Iub2z4 & Pub2z4);
assign Pub2z4 = (Wub2z4 & Dvb2z4);
assign Dvb2z4 = (Kvb2z4 & Xnjwx4);
assign Xnjwx4 = (~(Rvb2z4 & M66wx4));
assign Rvb2z4 = (~(J43wx4 | M3ovx4));
assign J43wx4 = (!Wdxvx4);
assign Kvb2z4 = (Una2z4 & Mn3wx4);
assign Una2z4 = (~(Yvb2z4 & Fwb2z4));
assign Yvb2z4 = (Ucqvx4 & O9qvx4);
assign Wub2z4 = (Zvyvx4 & Og4wx4);
assign Og4wx4 = (~(Mwb2z4 & Q5gvx4));
assign Mwb2z4 = (Huqvx4 & Kzxvx4);
assign Huqvx4 = (~(M3ovx4 | Us2wx4));
assign Zvyvx4 = (~(Twb2z4 & M66wx4));
assign M66wx4 = (Fjgvx4 & Z6gvx4);
assign Twb2z4 = (~(M3ovx4 | T93wx4));
assign Iub2z4 = (Axb2z4 & Hxb2z4);
assign Hxb2z4 = (Oxb2z4 & Yt3wx4);
assign Yt3wx4 = (~(Ucqvx4 & P6xvx4));
assign Oxb2z4 = (Vxb2z4 & Cyb2z4);
assign Cyb2z4 = (~(Mj8vx4 & Jyb2z4));
assign Jyb2z4 = (~(Qyb2z4 & Xyb2z4));
assign Xyb2z4 = (Ezb2z4 & Lzb2z4);
assign Lzb2z4 = (~(Nuewx4 & Szb2z4));
assign Szb2z4 = (S4xvx4 | Zzb2z4);
assign Nuewx4 = (~(Jhxvx4 | U9gvx4));
assign Ezb2z4 = (G0c2z4 & Xhiwx4);
assign Xhiwx4 = (~(N0c2z4 & Ju5wx4));
assign N0c2z4 = (~(S4xvx4 | Us2wx4));
assign G0c2z4 = (~(U0c2z4 & Ps3wx4));
assign U0c2z4 = (~(Cn8vx4 | Nggvx4));
assign Qyb2z4 = (B1c2z4 & I1c2z4);
assign I1c2z4 = (Pvewx4 | Gcqvx4);
assign B1c2z4 = (P1c2z4 & W1c2z4);
assign W1c2z4 = (~(A0zvx4 & D2c2z4));
assign D2c2z4 = (Nj4wx4 | K2c2z4);
assign K2c2z4 = (~(Msyvx4 | U9gvx4));
assign Msyvx4 = (R2c2z4 & Y2c2z4);
assign Y2c2z4 = (F3c2z4 & vis_pc_o[27]);
assign F3c2z4 = (Hx8vx4 & Rryvx4);
assign Rryvx4 = (~(Wgb2z4 & Rob2z4));
assign Rob2z4 = (Igb2z4 & Lzuvx4);
assign Lzuvx4 = (!vis_ipsr_o[3]);
assign Igb2z4 = (~(vis_ipsr_o[4] | vis_ipsr_o[5]));
assign Wgb2z4 = (Ckb2z4 & Xkuvx4);
assign Xkuvx4 = (!vis_ipsr_o[2]);
assign Ckb2z4 = (Gxqvx4 & T0rvx4);
assign T0rvx4 = (!vis_ipsr_o[1]);
assign Gxqvx4 = (!vis_ipsr_o[0]);
assign R2c2z4 = (M3c2z4 & vis_pc_o[30]);
assign M3c2z4 = (vis_pc_o[29] & vis_pc_o[28]);
assign P1c2z4 = (~(T3c2z4 & Zrvvx4));
assign T3c2z4 = (~(A4c2z4 & H4c2z4));
assign H4c2z4 = (~(C9yvx4 & O9qvx4));
assign A4c2z4 = (S87wx4 | F3ovx4);
assign Vxb2z4 = (~(O4c2z4 & Rexvx4));
assign Rexvx4 = (~(V4c2z4 | Fpmwx4));
assign Fpmwx4 = (!vis_pc_o[2]);
assign V4c2z4 = (~(Eg8vx4 & Efewx4));
assign Efewx4 = (!Ki8vx4);
assign O4c2z4 = (~(Pvewx4 | Gcqvx4));
assign Gcqvx4 = (!Fqlwx4);
assign Pvewx4 = (~(P9fwx4 & M3ovx4));
assign P9fwx4 = (P6xvx4 & Ujxvx4);
assign Axb2z4 = (C5c2z4 & J5c2z4);
assign J5c2z4 = (~(Eznvx4 & Kzxvx4));
assign C5c2z4 = (S4xvx4 ? X5c2z4 : Q5c2z4);
assign X5c2z4 = (E6c2z4 & L6c2z4);
assign L6c2z4 = (~(H0zvx4 & O9qvx4));
assign E6c2z4 = (S6c2z4 & Z6c2z4);
assign Z6c2z4 = (~(G7c2z4 & Q5gvx4));
assign G7c2z4 = (Wdqvx4 & Kzxvx4);
assign S6c2z4 = (~(R5dwx4 & P6xvx4));
assign Q5c2z4 = (R7qvx4 | T93wx4);
assign Bub2z4 = (Vlsvx4 ? U7c2z4 : N7c2z4);
assign Vlsvx4 = (!vis_pc_o[0]);
assign U7c2z4 = (Ipsvx4 & Zorvx4);
assign Zorvx4 = (!Hlsvx4);
assign Hlsvx4 = (A3gvx4 & B8c2z4);
assign N7c2z4 = (~(I8c2z4 & P8c2z4));
assign P8c2z4 = (~(Ipsvx4 & Wnnvx4));
assign Wnnvx4 = (~(I4gvx4 & B8c2z4));
assign B8c2z4 = (~(M9pvx4 & Dcrwx4));
assign M9pvx4 = (~(Kvfwx4 & W8c2z4));
assign W8c2z4 = (~(Qp3wx4 & B1ovx4));
assign Qp3wx4 = (U9gvx4 & Izwvx4);
assign Kvfwx4 = (N4yvx4 | Bl3wx4);
assign N4yvx4 = (!Howvx4);
assign Ipsvx4 = (~(Y8pvx4 & Dcrwx4));
assign Dcrwx4 = (~(D9c2z4 & K9c2z4));
assign K9c2z4 = (R9c2z4 & Y9c2z4);
assign Y9c2z4 = (Fac2z4 & Mac2z4);
assign Mac2z4 = (~(Tac2z4 & Abc2z4));
assign Abc2z4 = (~(Fpfwx4 | Bl3wx4));
assign Tac2z4 = (Wkxvx4 & Mj8vx4);
assign Wkxvx4 = (~(Efgvx4 | Whgvx4));
assign Fac2z4 = (Hbc2z4 & Gg7wx4);
assign Gg7wx4 = (~(Tlcwx4 & Xx2wx4));
assign Xx2wx4 = (U9gvx4 & U0ovx4);
assign Tlcwx4 = (~(Us2wx4 | Nggvx4));
assign Hbc2z4 = (~(Obc2z4 & Vbc2z4));
assign Vbc2z4 = (Hw2wx4 & W5yvx4);
assign Obc2z4 = (X77wx4 & Jwwvx4);
assign Jwwvx4 = (Mj8vx4 & F3ovx4);
assign R9c2z4 = (Ccc2z4 & Jcc2z4);
assign Jcc2z4 = (~(Qcc2z4 & R13wx4));
assign R13wx4 = (Rngwx4 & Z6gvx4);
assign Qcc2z4 = (Xcc2z4 & S87wx4);
assign Xcc2z4 = (Fqlwx4 | E44wx4);
assign E44wx4 = (~(Dbgvx4 | Efgvx4));
assign Fqlwx4 = (~(Dbgvx4 | Vdgvx4));
assign Ccc2z4 = (~(Edc2z4 & Z9dwx4));
assign Z9dwx4 = (~(Us2wx4 | Whgvx4));
assign Edc2z4 = (~(F3ovx4 | Fjgvx4));
assign D9c2z4 = (Ldc2z4 & Sdc2z4);
assign Sdc2z4 = (Zdc2z4 & Gec2z4);
assign Gec2z4 = (~(Nec2z4 & Pcyvx4));
assign Nec2z4 = (Nv6wx4 & Qx2wx4);
assign Zdc2z4 = (~(Rkgvx4 & Uec2z4));
assign Uec2z4 = (~(Wpsvx4 & Bfc2z4));
assign Bfc2z4 = (~(Ifc2z4 & O9qvx4));
assign Ifc2z4 = (~(M93wx4 | Db7wx4));
assign Db7wx4 = (!Ps3wx4);
assign Ps3wx4 = (~(B1ovx4 | Efgvx4));
assign Wpsvx4 = (Rkjwx4 & Pfc2z4);
assign Pfc2z4 = (~(Pxcwx4 & Trsvx4));
assign Pxcwx4 = (~(F3ovx4 | Bl3wx4));
assign Rkjwx4 = (Wt2wx4 | Hp2wx4);
assign Hp2wx4 = (!Trsvx4);
assign Trsvx4 = (~(R7qvx4 | Fjgvx4));
assign Ldc2z4 = (Wfc2z4 & Dgc2z4);
assign Dgc2z4 = (~(Y13wx4 & Kgc2z4));
assign Kgc2z4 = (~(Rgc2z4 & Ygc2z4));
assign Ygc2z4 = (~(Fhc2z4 | Whgvx4));
assign Rgc2z4 = (~(Nj4wx4 | Eznvx4));
assign Nj4wx4 = (~(B1ovx4 | Vdgvx4));
assign Y13wx4 = (~(Izwvx4 | Dmgvx4));
assign Wfc2z4 = (~(Vdgvx4 & Mhc2z4));
assign Mhc2z4 = (~(Thc2z4 & Aic2z4));
assign Aic2z4 = (Hic2z4 & Oic2z4);
assign Oic2z4 = (~(H0zvx4 | Zzfwx4));
assign Zzfwx4 = (~(Pxyvx4 | W5yvx4));
assign Pxyvx4 = (!P6xvx4);
assign Hic2z4 = (Vic2z4 & Cjc2z4);
assign Cjc2z4 = (~(Rkgvx4 & Jjc2z4));
assign Jjc2z4 = (~(Qjc2z4 & Xjc2z4));
assign Xjc2z4 = (~(Uj4wx4 & Rngwx4));
assign Uj4wx4 = (~(M93wx4 | Sh9vx4));
assign Qjc2z4 = (~(Ekc2z4 & F3ovx4));
assign Ekc2z4 = (~(Lkc2z4 & Skc2z4));
assign Skc2z4 = (~(Zkc2z4 & C2yvx4));
assign C2yvx4 = (O4ovx4 & Xmsvx4);
assign Xmsvx4 = (!Sh9vx4);
assign Zkc2z4 = (~(M3ovx4 | W7hwx4));
assign W7hwx4 = (Zn6wx4 & Glc2z4);
assign Glc2z4 = (C1svx4 | Ryrvx4);
assign Ryrvx4 = (!W49vx4);
assign C1svx4 = (!D69vx4);
assign Zn6wx4 = (~(N3svx4 | R89vx4));
assign N3svx4 = (!K79vx4);
assign Lkc2z4 = (~(Rngwx4 & Nlc2z4));
assign Nlc2z4 = (~(Ulc2z4 & Qqgwx4));
assign Qqgwx4 = (B8gwx4 & Bmc2z4);
assign Bmc2z4 = (Sh9vx4 | Aj9vx4);
assign B8gwx4 = (!O1jwx4);
assign O1jwx4 = (~(Bisvx4 | Sh9vx4));
assign Ulc2z4 = (Imc2z4 & H0kwx4);
assign H0kwx4 = (!Mgwvx4);
assign Mgwvx4 = (~(Ho8vx4 | Aj9vx4));
assign Imc2z4 = (~(Sh9vx4 & K8hwx4));
assign K8hwx4 = (Aj9vx4 & Bisvx4);
assign Bisvx4 = (!Cf9vx4);
assign Vic2z4 = (~(Wdqvx4 & Kzxvx4));
assign Wdqvx4 = (~(Mcgvx4 | Efgvx4));
assign Thc2z4 = (~(Pmc2z4 | Wmc2z4));
assign Wmc2z4 = (R7qvx4 ? Dnc2z4 : P6xvx4);
assign Dnc2z4 = (~(Wt2wx4 | B1ovx4));
assign Wt2wx4 = (!O9qvx4);
assign Pmc2z4 = (~(Knc2z4 & Rnc2z4));
assign Rnc2z4 = (Mvgwx4 | Mv2wx4);
assign Mv2wx4 = (!Zzb2z4);
assign Zzb2z4 = (~(Us2wx4 | Z6gvx4));
assign Knc2z4 = (~(B73wx4 & U9gvx4));
assign Y8pvx4 = (~(Keqvx4 & Ync2z4));
assign Ync2z4 = (~(P7pvx4 & Howvx4));
assign P7pvx4 = (~(Us2wx4 | U9gvx4));
assign I8c2z4 = (Izwvx4 | Xyfvx4);
assign Ema2z4 = (Oq42z4 | V3wvx4);
assign V3wvx4 = (!N5qvx4);
assign N5qvx4 = (~(Foc2z4 & Moc2z4));
assign Moc2z4 = (~(Gzvvx4 & Oxnvx4));
assign Oxnvx4 = (~(Toc2z4 & Apc2z4));
assign Apc2z4 = (~(Vb9wx4 & Hpc2z4));
assign Hpc2z4 = (~(Opc2z4 & Vpc2z4));
assign Vpc2z4 = (Cqc2z4 & Jqc2z4);
assign Jqc2z4 = (Qqc2z4 & Xqc2z4);
assign Xqc2z4 = (~(Zd9wx4 & vis_r14_o[0]));
assign Zd9wx4 = (~(Erc2z4 | Tja2z4));
assign Qqc2z4 = (~(Wf9wx4 & vis_r12_o[0]));
assign Wf9wx4 = (~(Lrc2z4 | Tja2z4));
assign Cqc2z4 = (Src2z4 & Zrc2z4);
assign Zrc2z4 = (~(Dg9wx4 & vis_r11_o[0]));
assign Dg9wx4 = (~(Gsc2z4 | Nsc2z4));
assign Src2z4 = (~(Mh9wx4 & vis_r10_o[0]));
assign Mh9wx4 = (~(Gsc2z4 | Erc2z4));
assign Opc2z4 = (Usc2z4 & Cawwx4);
assign Usc2z4 = (Btc2z4 & Itc2z4);
assign Itc2z4 = (~(Th9wx4 & vis_r9_o[0]));
assign Th9wx4 = (~(Gsc2z4 | Ptc2z4));
assign Btc2z4 = (~(Oi9wx4 & vis_r8_o[0]));
assign Oi9wx4 = (~(Gsc2z4 | Lrc2z4));
assign Gsc2z4 = (Wtc2z4 | Tjh2z4[2]);
assign Vb9wx4 = (Duc2z4 & Kuc2z4);
assign Toc2z4 = (~(Qj9wx4 & Kycvx4));
assign Qj9wx4 = (~(Jj9wx4 | Kuc2z4));
assign Kuc2z4 = (Ruc2z4 & Yuc2z4);
assign Yuc2z4 = (~(Fvc2z4 | Huiwx4));
assign Huiwx4 = (~(M93wx4 | Zrvvx4));
assign Fvc2z4 = (~(Mvc2z4 & Keqvx4));
assign Keqvx4 = (!Xkfwx4);
assign Xkfwx4 = (~(Tv2wx4 | Zrvvx4));
assign Tv2wx4 = (!X43wx4);
assign X43wx4 = (~(S4xvx4 | U9gvx4));
assign Mvc2z4 = (Nsc2z4 | Tja2z4);
assign Tja2z4 = (~(Tjh2z4[3] & Tjh2z4[2]));
assign Ruc2z4 = (Tvc2z4 & Awc2z4);
assign Awc2z4 = (Bl3wx4 ? Owc2z4 : Hwc2z4);
assign Owc2z4 = (~(Ffqvx4 & M3ovx4));
assign Ffqvx4 = (Ucqvx4 & F3ovx4);
assign Ucqvx4 = (Nggvx4 & S4xvx4);
assign Hwc2z4 = (Xviwx4 | Vdgvx4);
assign Xviwx4 = (!Eiqvx4);
assign Eiqvx4 = (~(Zj3wx4 | Mcgvx4));
assign Tvc2z4 = (Vwc2z4 & Cxc2z4);
assign Cxc2z4 = (~(Jxc2z4 & Ncqvx4));
assign Jxc2z4 = (~(Fpfwx4 | Cn8vx4));
assign Vwc2z4 = (~(B1ovx4 & Qxc2z4));
assign Qxc2z4 = (P6xvx4 | O9qvx4);
assign P6xvx4 = (~(Zrvvx4 | Z6gvx4));
assign Jj9wx4 = (!Duc2z4);
assign Gzvvx4 = (Xxc2z4 & D7qvx4);
assign Xxc2z4 = (~(Eyc2z4 & Lyc2z4));
assign Lyc2z4 = (Syc2z4 & Zyc2z4);
assign Zyc2z4 = (~(Gzc2z4 & F3ovx4));
assign Gzc2z4 = (~(Q68wx4 & Nzc2z4));
assign Nzc2z4 = (Oedwx4 | H33wx4);
assign H33wx4 = (!Wxcwx4);
assign Wxcwx4 = (~(B1ovx4 | Mcgvx4));
assign Oedwx4 = (!Eznvx4);
assign Eznvx4 = (~(Bl3wx4 | Efgvx4));
assign Q68wx4 = (!Ujiwx4);
assign Ujiwx4 = (~(M93wx4 | Dbgvx4));
assign Syc2z4 = (Uzc2z4 & Tscwx4);
assign Tscwx4 = (B0d2z4 | Duc2z4);
assign B0d2z4 = (!I0d2z4);
assign Uzc2z4 = (~(P0d2z4 & I7pvx4));
assign I7pvx4 = (~(F3ovx4 | U9gvx4));
assign P0d2z4 = (~(Mcgvx4 | Fjgvx4));
assign Eyc2z4 = (W0d2z4 & D1d2z4);
assign D1d2z4 = (~(H0zvx4 & S4xvx4));
assign W0d2z4 = (K1d2z4 & R1d2z4);
assign R1d2z4 = (Acfwx4 | Efgvx4);
assign Acfwx4 = (!Uvrwx4);
assign Uvrwx4 = (~(M3ovx4 | Zrvvx4));
assign K1d2z4 = (~(Jp3wx4 & U9gvx4));
assign Jp3wx4 = (B1vvx4 & Dbgvx4);
assign Foc2z4 = (~(Dmh2z4[0] & K1wvx4));
assign K1wvx4 = (Y1d2z4 & D7qvx4);
assign D7qvx4 = (!Mrsvx4);
assign Mrsvx4 = (F2d2z4 & M2d2z4);
assign M2d2z4 = (T2d2z4 & A3d2z4);
assign A3d2z4 = (H3d2z4 & O3d2z4);
assign O3d2z4 = (~(V3d2z4 & P5yvx4));
assign P5yvx4 = (~(S4xvx4 | Zrvvx4));
assign V3d2z4 = (~(Dmgvx4 | Nggvx4));
assign H3d2z4 = (C4d2z4 & Mn3wx4);
assign C4d2z4 = (~(Whgvx4 & J4d2z4));
assign J4d2z4 = (Q4d2z4 | Zmewx4);
assign Zmewx4 = (C9yvx4 & Xhqvx4);
assign C9yvx4 = (X4d2z4 & Izwvx4);
assign X4d2z4 = (~(Mcgvx4 | Vdgvx4));
assign Q4d2z4 = (Vdgvx4 ? H0zvx4 : Xfkwx4);
assign H0zvx4 = (~(Zj3wx4 | M93wx4));
assign Zj3wx4 = (!Sy2wx4);
assign Sy2wx4 = (~(Us2wx4 | Dbgvx4));
assign Xfkwx4 = (Ju5wx4 & Hgxvx4);
assign Hgxvx4 = (!Q5gvx4);
assign T2d2z4 = (E5d2z4 & L5d2z4);
assign L5d2z4 = (~(S5d2z4 & Howvx4));
assign Howvx4 = (~(S4xvx4 | Cn8vx4));
assign S5d2z4 = (~(B1ovx4 | Z6gvx4));
assign E5d2z4 = (Z5d2z4 & G6d2z4);
assign G6d2z4 = (~(N6d2z4 & Pkxvx4));
assign N6d2z4 = (~(S87wx4 | Mj8vx4));
assign Z5d2z4 = (~(U6d2z4 & Fwb2z4));
assign Fwb2z4 = (~(M93wx4 | Efgvx4));
assign U6d2z4 = (~(Jhxvx4 | Sr2wx4));
assign Sr2wx4 = (!Qx2wx4);
assign Qx2wx4 = (B1ovx4 & W5yvx4);
assign F2d2z4 = (B7d2z4 & I7d2z4);
assign I7d2z4 = (Ru52z4 & P7d2z4);
assign P7d2z4 = (~(W7d2z4 & D8d2z4));
assign D8d2z4 = (~(T93wx4 | Vdgvx4));
assign W7d2z4 = (Mcgvx4 & Ju5wx4);
assign Ju5wx4 = (Kzxvx4 & Z6gvx4);
assign Kzxvx4 = (Fjgvx4 & Nggvx4);
assign Ru52z4 = (~(Aq1wx4 | Ry5wx4));
assign Ry5wx4 = (Jtkwx4 & Clewx4);
assign Clewx4 = (!Jppvx4);
assign Jppvx4 = (~(B73wx4 & Izwvx4));
assign B73wx4 = (Dbgvx4 & O4ovx4);
assign Jtkwx4 = (~(Efgvx4 | Nggvx4));
assign Aq1wx4 = (~(Hq1wx4 | F3ovx4));
assign Hq1wx4 = (!B1vvx4);
assign B1vvx4 = (~(Mcgvx4 | Nggvx4));
assign B7d2z4 = (K8d2z4 & Ol6wx4);
assign Ol6wx4 = (R8d2z4 & Lbiwx4);
assign Lbiwx4 = (Zrvvx4 | B1ovx4);
assign R8d2z4 = (~(Ncqvx4 & Y8d2z4));
assign Y8d2z4 = (I3swx4 | T1xvx4);
assign T1xvx4 = (~(Sznvx4 | F3ovx4));
assign I3swx4 = (~(Ujxvx4 | Sznvx4));
assign Sznvx4 = (!Pkxvx4);
assign Pkxvx4 = (~(Zrvvx4 | Vdgvx4));
assign Ujxvx4 = (!Fjewx4);
assign Fjewx4 = (F9d2z4 & M9d2z4);
assign M9d2z4 = (T9d2z4 & Aad2z4);
assign Aad2z4 = (~(Azrwx4 | Ilwvx4));
assign Ilwvx4 = (~(B5cwx4 | G6wvx4));
assign G6wvx4 = (!Ot9vx4);
assign Azrwx4 = (Ks9vx4 & Q0lwx4);
assign Q0lwx4 = (X9yvx4 | Gr9vx4);
assign T9d2z4 = (~(Qtrwx4 | Dxrwx4));
assign Dxrwx4 = (Gr9vx4 & X9yvx4);
assign X9yvx4 = (~(X0lwx4 & Cwawx4));
assign Qtrwx4 = (~(Cwawx4 | X0lwx4));
assign X0lwx4 = (~(S1lwx4 | Yo9vx4));
assign Cwawx4 = (!Cq9vx4);
assign F9d2z4 = (Had2z4 & Oad2z4);
assign Oad2z4 = (~(Su9vx4 & Vad2z4));
assign Vad2z4 = (Wv9vx4 | Ot9vx4);
assign Had2z4 = (~(E4xvx4 | Vklwx4));
assign Vklwx4 = (~(Xy8wx4 | Layvx4));
assign Layvx4 = (!S1lwx4);
assign S1lwx4 = (~(Sayvx4 & Dmwvx4));
assign E4xvx4 = (~(Dmwvx4 | Sayvx4));
assign Sayvx4 = (Cbd2z4 & B5cwx4);
assign B5cwx4 = (!Wv9vx4);
assign Cbd2z4 = (~(Ot9vx4 | Su9vx4));
assign Dmwvx4 = (!Bx9vx4);
assign K8d2z4 = (Jbd2z4 & Qbd2z4);
assign Qbd2z4 = (~(Xbd2z4 & A0zvx4));
assign A0zvx4 = (~(Jhxvx4 | F3ovx4));
assign Jhxvx4 = (!Z7fwx4);
assign Z7fwx4 = (~(Cn8vx4 | Fjgvx4));
assign Xbd2z4 = (~(Mvgwx4 | Bl3wx4));
assign Mvgwx4 = (!Qaqvx4);
assign Qaqvx4 = (~(Mj8vx4 | Dmgvx4));
assign Jbd2z4 = (~(O76wx4 & P03wx4));
assign O76wx4 = (Xhqvx4 & Izwvx4);
assign Xhqvx4 = (Rngwx4 & R7qvx4);
assign R7qvx4 = (!Dmgvx4);
assign Rngwx4 = (O4ovx4 & Zrvvx4);
assign O4ovx4 = (!Mj8vx4);
assign Y1d2z4 = (~(Ecd2z4 & Lcd2z4));
assign Lcd2z4 = (Scd2z4 & Zcd2z4);
assign Zcd2z4 = (Gdd2z4 & Ndd2z4);
assign Ndd2z4 = (~(Hrewx4 & Nv6wx4));
assign Nv6wx4 = (Us2wx4 & Zrvvx4);
assign Zrvvx4 = (!Fjgvx4);
assign Hrewx4 = (~(M3ovx4 | Vdgvx4));
assign M3ovx4 = (!Mcgvx4);
assign Gdd2z4 = (~(Ax0xx4 | Wdxvx4));
assign Wdxvx4 = (~(U9gvx4 | Nggvx4));
assign Ax0xx4 = (~(Dbgvx4 | Mcgvx4));
assign Scd2z4 = (L9dwx4 & Udd2z4);
assign Udd2z4 = (~(Z6gvx4 & Bed2z4));
assign Bed2z4 = (Vdgvx4 | Zocwx4);
assign Zocwx4 = (~(Bl3wx4 | B1ovx4));
assign L9dwx4 = (Ph7wx4 | U9gvx4);
assign Ph7wx4 = (!H5mwx4);
assign Ecd2z4 = (Ied2z4 & Ped2z4);
assign Ped2z4 = (Wed2z4 & Omcwx4);
assign Omcwx4 = (I0d2z4 | Duc2z4);
assign Duc2z4 = (Dfd2z4 & Kfd2z4);
assign Kfd2z4 = (~(Rfd2z4 & P03wx4));
assign P03wx4 = (Bl3wx4 & S4xvx4);
assign S4xvx4 = (!Vdgvx4);
assign Bl3wx4 = (!U9gvx4);
assign Rfd2z4 = (Cn8vx4 & Hw2wx4);
assign Dfd2z4 = (Mn3wx4 | Mj8vx4);
assign Mn3wx4 = (~(V6swx4 & Pcyvx4));
assign Pcyvx4 = (Mcgvx4 & Izwvx4);
assign Izwvx4 = (!Cn8vx4);
assign V6swx4 = (Yfd2z4 & O9qvx4);
assign O9qvx4 = (~(U0ovx4 | Z6gvx4));
assign Yfd2z4 = (~(E78wx4 | Us2wx4));
assign I0d2z4 = (Xy8wx4 ? Mgd2z4 : Fgd2z4);
assign Xy8wx4 = (!Yo9vx4);
assign Mgd2z4 = (Un9vx4 ? Ahd2z4 : Tgd2z4);
assign Ahd2z4 = (Yryvx4 ? Ohd2z4 : Hhd2z4);
assign Ohd2z4 = (Vhd2z4 & Cid2z4);
assign Cid2z4 = (Jid2z4 & Qid2z4);
assign Qid2z4 = (~(H9xvx4 & Rzpwx4));
assign Rzpwx4 = (!D9uwx4);
assign D9uwx4 = (Xid2z4 & Ejd2z4);
assign Ejd2z4 = (Ljd2z4 & Sjd2z4);
assign Sjd2z4 = (Zjd2z4 & Gkd2z4);
assign Gkd2z4 = (~(Nkd2z4 & vis_r2_o[21]));
assign Zjd2z4 = (~(Ukd2z4 & vis_r6_o[21]));
assign Ljd2z4 = (Bld2z4 & Ild2z4);
assign Ild2z4 = (~(Pld2z4 & vis_r5_o[21]));
assign Bld2z4 = (~(Wld2z4 & vis_r4_o[21]));
assign Xid2z4 = (Dmd2z4 & Kmd2z4);
assign Kmd2z4 = (Rmd2z4 & Ymd2z4);
assign Ymd2z4 = (~(Fnd2z4 & vis_r1_o[21]));
assign Rmd2z4 = (~(Mnd2z4 & vis_r0_o[21]));
assign Dmd2z4 = (Tnd2z4 & Aod2z4);
assign Aod2z4 = (~(Hod2z4 & vis_r3_o[21]));
assign Tnd2z4 = (~(Ood2z4 & vis_r7_o[21]));
assign Jid2z4 = (~(Spqvx4 & Y9uwx4));
assign Y9uwx4 = (!G4qwx4);
assign G4qwx4 = (Vod2z4 & Cpd2z4);
assign Cpd2z4 = (Jpd2z4 & Qpd2z4);
assign Qpd2z4 = (Xpd2z4 & Eqd2z4);
assign Eqd2z4 = (~(Nkd2z4 & vis_r2_o[22]));
assign Xpd2z4 = (~(Ukd2z4 & vis_r6_o[22]));
assign Jpd2z4 = (Lqd2z4 & Sqd2z4);
assign Sqd2z4 = (~(Pld2z4 & vis_r5_o[22]));
assign Lqd2z4 = (~(Wld2z4 & vis_r4_o[22]));
assign Vod2z4 = (Zqd2z4 & Grd2z4);
assign Grd2z4 = (Nrd2z4 & Urd2z4);
assign Urd2z4 = (~(Fnd2z4 & vis_r1_o[22]));
assign Nrd2z4 = (~(Mnd2z4 & vis_r0_o[22]));
assign Zqd2z4 = (Bsd2z4 & Isd2z4);
assign Isd2z4 = (~(Hod2z4 & vis_r3_o[22]));
assign Bsd2z4 = (~(Ood2z4 & vis_r7_o[22]));
assign Vhd2z4 = (Psd2z4 & Wsd2z4);
assign Wsd2z4 = (~(Lpqvx4 & N4qwx4));
assign N4qwx4 = (!Icxwx4);
assign Icxwx4 = (Dtd2z4 & Ktd2z4);
assign Ktd2z4 = (Rtd2z4 & Ytd2z4);
assign Ytd2z4 = (Fud2z4 & Mud2z4);
assign Mud2z4 = (~(vis_r2_o[23] & Nkd2z4));
assign Fud2z4 = (~(vis_r6_o[23] & Ukd2z4));
assign Rtd2z4 = (Tud2z4 & Avd2z4);
assign Avd2z4 = (~(vis_r5_o[23] & Pld2z4));
assign Tud2z4 = (~(vis_r4_o[23] & Wld2z4));
assign Dtd2z4 = (Hvd2z4 & Ovd2z4);
assign Ovd2z4 = (Vvd2z4 & Cwd2z4);
assign Cwd2z4 = (~(vis_r1_o[23] & Fnd2z4));
assign Vvd2z4 = (~(vis_r0_o[23] & Mnd2z4));
assign Hvd2z4 = (Jwd2z4 & Qwd2z4);
assign Qwd2z4 = (~(vis_r3_o[23] & Hod2z4));
assign Jwd2z4 = (~(vis_r7_o[23] & Ood2z4));
assign Psd2z4 = (~(Onwwx4 & L3qwx4));
assign L3qwx4 = (!Mnvwx4);
assign Mnvwx4 = (Xwd2z4 & Exd2z4);
assign Exd2z4 = (Lxd2z4 & Sxd2z4);
assign Sxd2z4 = (Zxd2z4 & Gyd2z4);
assign Gyd2z4 = (~(vis_r2_o[24] & Nkd2z4));
assign Zxd2z4 = (~(vis_r6_o[24] & Ukd2z4));
assign Lxd2z4 = (Nyd2z4 & Uyd2z4);
assign Uyd2z4 = (~(vis_r5_o[24] & Pld2z4));
assign Nyd2z4 = (~(vis_r4_o[24] & Wld2z4));
assign Xwd2z4 = (Bzd2z4 & Izd2z4);
assign Izd2z4 = (Pzd2z4 & Wzd2z4);
assign Wzd2z4 = (~(vis_r1_o[24] & Fnd2z4));
assign Pzd2z4 = (~(vis_r0_o[24] & Mnd2z4));
assign Bzd2z4 = (D0e2z4 & K0e2z4);
assign K0e2z4 = (~(vis_r3_o[24] & Hod2z4));
assign D0e2z4 = (~(vis_r7_o[24] & Ood2z4));
assign Hhd2z4 = (R0e2z4 & Y0e2z4);
assign Y0e2z4 = (F1e2z4 & M1e2z4);
assign M1e2z4 = (~(H9xvx4 & Flqwx4));
assign Flqwx4 = (!Xcuwx4);
assign Xcuwx4 = (T1e2z4 & A2e2z4);
assign A2e2z4 = (H2e2z4 & O2e2z4);
assign O2e2z4 = (V2e2z4 & C3e2z4);
assign C3e2z4 = (~(Nkd2z4 & vis_r2_o[17]));
assign V2e2z4 = (~(Ukd2z4 & vis_r6_o[17]));
assign H2e2z4 = (J3e2z4 & Q3e2z4);
assign Q3e2z4 = (~(Pld2z4 & vis_r5_o[17]));
assign J3e2z4 = (~(Wld2z4 & vis_r4_o[17]));
assign T1e2z4 = (X3e2z4 & E4e2z4);
assign E4e2z4 = (L4e2z4 & S4e2z4);
assign S4e2z4 = (~(Fnd2z4 & vis_r1_o[17]));
assign L4e2z4 = (~(Mnd2z4 & vis_r0_o[17]));
assign X3e2z4 = (Z4e2z4 & G5e2z4);
assign G5e2z4 = (~(Hod2z4 & vis_r3_o[17]));
assign Z4e2z4 = (~(Ood2z4 & vis_r7_o[17]));
assign F1e2z4 = (~(Spqvx4 & Sduwx4));
assign Sduwx4 = (!H1qwx4);
assign H1qwx4 = (N5e2z4 & U5e2z4);
assign U5e2z4 = (B6e2z4 & I6e2z4);
assign I6e2z4 = (P6e2z4 & W6e2z4);
assign W6e2z4 = (~(Nkd2z4 & vis_r2_o[18]));
assign P6e2z4 = (~(Ukd2z4 & vis_r6_o[18]));
assign B6e2z4 = (D7e2z4 & K7e2z4);
assign K7e2z4 = (~(Pld2z4 & vis_r5_o[18]));
assign D7e2z4 = (~(Wld2z4 & vis_r4_o[18]));
assign N5e2z4 = (R7e2z4 & Y7e2z4);
assign Y7e2z4 = (F8e2z4 & M8e2z4);
assign M8e2z4 = (~(Fnd2z4 & vis_r1_o[18]));
assign F8e2z4 = (~(Mnd2z4 & vis_r0_o[18]));
assign R7e2z4 = (T8e2z4 & A9e2z4);
assign A9e2z4 = (~(Hod2z4 & vis_r3_o[18]));
assign T8e2z4 = (~(Ood2z4 & vis_r7_o[18]));
assign R0e2z4 = (H9e2z4 & O9e2z4);
assign O9e2z4 = (~(Lpqvx4 & F0qwx4));
assign F0qwx4 = (!Bjxwx4);
assign Bjxwx4 = (V9e2z4 & Cae2z4);
assign Cae2z4 = (Jae2z4 & Qae2z4);
assign Qae2z4 = (Xae2z4 & Ebe2z4);
assign Ebe2z4 = (~(Nkd2z4 & vis_r2_o[19]));
assign Xae2z4 = (~(Ukd2z4 & vis_r6_o[19]));
assign Jae2z4 = (Lbe2z4 & Sbe2z4);
assign Sbe2z4 = (~(Pld2z4 & vis_r5_o[19]));
assign Lbe2z4 = (~(Wld2z4 & vis_r4_o[19]));
assign V9e2z4 = (Zbe2z4 & Gce2z4);
assign Gce2z4 = (Nce2z4 & Uce2z4);
assign Uce2z4 = (~(Fnd2z4 & vis_r1_o[19]));
assign Nce2z4 = (~(Mnd2z4 & vis_r0_o[19]));
assign Zbe2z4 = (Bde2z4 & Ide2z4);
assign Ide2z4 = (~(Hod2z4 & vis_r3_o[19]));
assign Bde2z4 = (~(Ood2z4 & vis_r7_o[19]));
assign H9e2z4 = (~(Onwwx4 & V1qwx4));
assign V1qwx4 = (!Dmvwx4);
assign Dmvwx4 = (Pde2z4 & Wde2z4);
assign Wde2z4 = (Dee2z4 & Kee2z4);
assign Kee2z4 = (Ree2z4 & Yee2z4);
assign Yee2z4 = (~(Nkd2z4 & vis_r2_o[20]));
assign Ree2z4 = (~(Ukd2z4 & vis_r6_o[20]));
assign Dee2z4 = (Ffe2z4 & Mfe2z4);
assign Mfe2z4 = (~(Pld2z4 & vis_r5_o[20]));
assign Ffe2z4 = (~(Wld2z4 & vis_r4_o[20]));
assign Pde2z4 = (Tfe2z4 & Age2z4);
assign Age2z4 = (Hge2z4 & Oge2z4);
assign Oge2z4 = (~(Fnd2z4 & vis_r1_o[20]));
assign Hge2z4 = (~(Mnd2z4 & vis_r0_o[20]));
assign Tfe2z4 = (Vge2z4 & Che2z4);
assign Che2z4 = (~(Hod2z4 & vis_r3_o[20]));
assign Vge2z4 = (~(Ood2z4 & vis_r7_o[20]));
assign Tgd2z4 = (Yryvx4 ? Qhe2z4 : Jhe2z4);
assign Qhe2z4 = (Xhe2z4 & Eie2z4);
assign Eie2z4 = (Lie2z4 & Sie2z4);
assign Sie2z4 = (~(H9xvx4 & Ddqwx4));
assign Ddqwx4 = (!Eruwx4);
assign Eruwx4 = (Zie2z4 & Gje2z4);
assign Gje2z4 = (Nje2z4 & Uje2z4);
assign Uje2z4 = (Bke2z4 & Ike2z4);
assign Ike2z4 = (~(vis_r2_o[29] & Nkd2z4));
assign Bke2z4 = (~(vis_r6_o[29] & Ukd2z4));
assign Nje2z4 = (Pke2z4 & Wke2z4);
assign Wke2z4 = (~(vis_r5_o[29] & Pld2z4));
assign Pke2z4 = (~(vis_r4_o[29] & Wld2z4));
assign Zie2z4 = (Dle2z4 & Kle2z4);
assign Kle2z4 = (Rle2z4 & Yle2z4);
assign Yle2z4 = (~(vis_r1_o[29] & Fnd2z4));
assign Rle2z4 = (~(vis_r0_o[29] & Mnd2z4));
assign Dle2z4 = (Fme2z4 & Mme2z4);
assign Mme2z4 = (~(vis_r3_o[29] & Hod2z4));
assign Fme2z4 = (~(vis_r7_o[29] & Ood2z4));
assign Lie2z4 = (~(Spqvx4 & Zruwx4));
assign Zruwx4 = (!Saqwx4);
assign Saqwx4 = (Tme2z4 & Ane2z4);
assign Ane2z4 = (Hne2z4 & One2z4);
assign One2z4 = (Vne2z4 & Coe2z4);
assign Coe2z4 = (~(vis_r2_o[30] & Nkd2z4));
assign Vne2z4 = (~(vis_r6_o[30] & Ukd2z4));
assign Hne2z4 = (Joe2z4 & Qoe2z4);
assign Qoe2z4 = (~(vis_r5_o[30] & Pld2z4));
assign Joe2z4 = (~(vis_r4_o[30] & Wld2z4));
assign Tme2z4 = (Xoe2z4 & Epe2z4);
assign Epe2z4 = (Lpe2z4 & Spe2z4);
assign Spe2z4 = (~(vis_r1_o[30] & Fnd2z4));
assign Lpe2z4 = (~(vis_r0_o[30] & Mnd2z4));
assign Xoe2z4 = (Zpe2z4 & Gqe2z4);
assign Gqe2z4 = (~(vis_r3_o[30] & Hod2z4));
assign Zpe2z4 = (~(vis_r7_o[30] & Ood2z4));
assign Xhe2z4 = (Nqe2z4 & Uqe2z4);
assign Uqe2z4 = (~(Lpqvx4 & Nbqwx4));
assign Nbqwx4 = (!N3ywx4);
assign N3ywx4 = (Bre2z4 & Ire2z4);
assign Ire2z4 = (Pre2z4 & Wre2z4);
assign Wre2z4 = (Dse2z4 & Kse2z4);
assign Kse2z4 = (~(Nkd2z4 & vis_r2_o[31]));
assign Dse2z4 = (~(Ukd2z4 & vis_r6_o[31]));
assign Pre2z4 = (Rse2z4 & Yse2z4);
assign Yse2z4 = (~(Pld2z4 & vis_r5_o[31]));
assign Rse2z4 = (~(Wld2z4 & vis_r4_o[31]));
assign Bre2z4 = (Fte2z4 & Mte2z4);
assign Mte2z4 = (Tte2z4 & Aue2z4);
assign Aue2z4 = (~(Fnd2z4 & vis_r1_o[31]));
assign Tte2z4 = (~(Mnd2z4 & vis_r0_o[31]));
assign Fte2z4 = (Hue2z4 & Oue2z4);
assign Oue2z4 = (~(Hod2z4 & vis_r3_o[31]));
assign Hue2z4 = (~(Ood2z4 & vis_r7_o[31]));
assign Nqe2z4 = (~(Onwwx4 & Laqwx4));
assign Laqwx4 = (!Cawwx4);
assign Cawwx4 = (Vue2z4 & Cve2z4);
assign Cve2z4 = (Jve2z4 & Qve2z4);
assign Qve2z4 = (Xve2z4 & Ewe2z4);
assign Ewe2z4 = (~(Nkd2z4 & vis_r2_o[0]));
assign Xve2z4 = (~(Ukd2z4 & vis_r6_o[0]));
assign Jve2z4 = (Lwe2z4 & Swe2z4);
assign Swe2z4 = (~(Pld2z4 & vis_r5_o[0]));
assign Lwe2z4 = (~(Wld2z4 & vis_r4_o[0]));
assign Vue2z4 = (Zwe2z4 & Gxe2z4);
assign Gxe2z4 = (Nxe2z4 & Uxe2z4);
assign Uxe2z4 = (~(Fnd2z4 & vis_r1_o[0]));
assign Nxe2z4 = (~(Mnd2z4 & vis_r0_o[0]));
assign Zwe2z4 = (Bye2z4 & Iye2z4);
assign Iye2z4 = (~(Hod2z4 & vis_r3_o[0]));
assign Bye2z4 = (~(Ood2z4 & vis_r7_o[0]));
assign Jhe2z4 = (Pye2z4 & Wye2z4);
assign Wye2z4 = (Dze2z4 & Kze2z4);
assign Kze2z4 = (~(H9xvx4 & E3qwx4));
assign E3qwx4 = (!U7uwx4);
assign U7uwx4 = (Rze2z4 & Yze2z4);
assign Yze2z4 = (F0f2z4 & M0f2z4);
assign M0f2z4 = (T0f2z4 & A1f2z4);
assign A1f2z4 = (~(Nkd2z4 & vis_r2_o[25]));
assign T0f2z4 = (~(Ukd2z4 & vis_r6_o[25]));
assign F0f2z4 = (H1f2z4 & O1f2z4);
assign O1f2z4 = (~(Pld2z4 & vis_r5_o[25]));
assign H1f2z4 = (~(Wld2z4 & vis_r4_o[25]));
assign Rze2z4 = (V1f2z4 & C2f2z4);
assign C2f2z4 = (J2f2z4 & Q2f2z4);
assign Q2f2z4 = (~(Fnd2z4 & vis_r1_o[25]));
assign J2f2z4 = (~(Mnd2z4 & vis_r0_o[25]));
assign V1f2z4 = (X2f2z4 & E3f2z4);
assign E3f2z4 = (~(Hod2z4 & vis_r3_o[25]));
assign X2f2z4 = (~(Ood2z4 & vis_r7_o[25]));
assign Dze2z4 = (~(Spqvx4 & Z6uwx4));
assign Z6uwx4 = (!Feqwx4);
assign Feqwx4 = (L3f2z4 & S3f2z4);
assign S3f2z4 = (Z3f2z4 & G4f2z4);
assign G4f2z4 = (N4f2z4 & U4f2z4);
assign U4f2z4 = (~(Nkd2z4 & vis_r2_o[26]));
assign N4f2z4 = (~(Ukd2z4 & vis_r6_o[26]));
assign Z3f2z4 = (B5f2z4 & I5f2z4);
assign I5f2z4 = (~(Pld2z4 & vis_r5_o[26]));
assign B5f2z4 = (~(Wld2z4 & vis_r4_o[26]));
assign L3f2z4 = (P5f2z4 & W5f2z4);
assign W5f2z4 = (D6f2z4 & K6f2z4);
assign K6f2z4 = (~(Fnd2z4 & vis_r1_o[26]));
assign D6f2z4 = (~(Mnd2z4 & vis_r0_o[26]));
assign P5f2z4 = (R6f2z4 & Y6f2z4);
assign Y6f2z4 = (~(Hod2z4 & vis_r3_o[26]));
assign R6f2z4 = (~(Ood2z4 & vis_r7_o[26]));
assign Pye2z4 = (F7f2z4 & M7f2z4);
assign M7f2z4 = (~(Lpqvx4 & Kdqwx4));
assign Kdqwx4 = (!Fexwx4);
assign Fexwx4 = (T7f2z4 & A8f2z4);
assign A8f2z4 = (H8f2z4 & O8f2z4);
assign O8f2z4 = (V8f2z4 & C9f2z4);
assign C9f2z4 = (~(vis_r2_o[27] & Nkd2z4));
assign V8f2z4 = (~(vis_r6_o[27] & Ukd2z4));
assign H8f2z4 = (J9f2z4 & Q9f2z4);
assign Q9f2z4 = (~(vis_r5_o[27] & Pld2z4));
assign J9f2z4 = (~(vis_r4_o[27] & Wld2z4));
assign T7f2z4 = (X9f2z4 & Eaf2z4);
assign Eaf2z4 = (Laf2z4 & Saf2z4);
assign Saf2z4 = (~(vis_r1_o[27] & Fnd2z4));
assign Laf2z4 = (~(vis_r0_o[27] & Mnd2z4));
assign X9f2z4 = (Zaf2z4 & Gbf2z4);
assign Gbf2z4 = (~(vis_r3_o[27] & Hod2z4));
assign Zaf2z4 = (~(vis_r7_o[27] & Ood2z4));
assign F7f2z4 = (~(Onwwx4 & Meqwx4));
assign Meqwx4 = (!F8wwx4);
assign F8wwx4 = (Nbf2z4 & Ubf2z4);
assign Ubf2z4 = (Bcf2z4 & Icf2z4);
assign Icf2z4 = (Pcf2z4 & Wcf2z4);
assign Wcf2z4 = (~(vis_r2_o[28] & Nkd2z4));
assign Pcf2z4 = (~(vis_r6_o[28] & Ukd2z4));
assign Bcf2z4 = (Ddf2z4 & Kdf2z4);
assign Kdf2z4 = (~(vis_r5_o[28] & Pld2z4));
assign Ddf2z4 = (~(vis_r4_o[28] & Wld2z4));
assign Nbf2z4 = (Rdf2z4 & Ydf2z4);
assign Ydf2z4 = (Fef2z4 & Mef2z4);
assign Mef2z4 = (~(vis_r1_o[28] & Fnd2z4));
assign Fef2z4 = (~(vis_r0_o[28] & Mnd2z4));
assign Rdf2z4 = (Tef2z4 & Aff2z4);
assign Aff2z4 = (~(vis_r3_o[28] & Hod2z4));
assign Tef2z4 = (~(vis_r7_o[28] & Ood2z4));
assign Fgd2z4 = (Un9vx4 ? Off2z4 : Hff2z4);
assign Off2z4 = (Yryvx4 ? Cgf2z4 : Vff2z4);
assign Cgf2z4 = (Jgf2z4 & Qgf2z4);
assign Qgf2z4 = (Xgf2z4 & Ehf2z4);
assign Ehf2z4 = (~(H9xvx4 & Bqqwx4));
assign Bqqwx4 = (!Qxuwx4);
assign Qxuwx4 = (Lhf2z4 & Shf2z4);
assign Shf2z4 = (Zhf2z4 & Gif2z4);
assign Gif2z4 = (Nif2z4 & Uif2z4);
assign Uif2z4 = (~(vis_r2_o[5] & Nkd2z4));
assign Nif2z4 = (~(vis_r6_o[5] & Ukd2z4));
assign Zhf2z4 = (Bjf2z4 & Ijf2z4);
assign Ijf2z4 = (~(vis_r5_o[5] & Pld2z4));
assign Bjf2z4 = (~(vis_r4_o[5] & Wld2z4));
assign Lhf2z4 = (Pjf2z4 & Wjf2z4);
assign Wjf2z4 = (Dkf2z4 & Kkf2z4);
assign Kkf2z4 = (~(vis_r1_o[5] & Fnd2z4));
assign Dkf2z4 = (~(vis_r0_o[5] & Mnd2z4));
assign Pjf2z4 = (Rkf2z4 & Ykf2z4);
assign Ykf2z4 = (~(vis_r3_o[5] & Hod2z4));
assign Rkf2z4 = (~(vis_r7_o[5] & Ood2z4));
assign Xgf2z4 = (~(Spqvx4 & Lyuwx4));
assign Lyuwx4 = (!Svqwx4);
assign Svqwx4 = (Flf2z4 & Mlf2z4);
assign Mlf2z4 = (Tlf2z4 & Amf2z4);
assign Amf2z4 = (Hmf2z4 & Omf2z4);
assign Omf2z4 = (~(Nkd2z4 & vis_r2_o[6]));
assign Hmf2z4 = (~(Ukd2z4 & vis_r6_o[6]));
assign Tlf2z4 = (Vmf2z4 & Cnf2z4);
assign Cnf2z4 = (~(Pld2z4 & vis_r5_o[6]));
assign Vmf2z4 = (~(Wld2z4 & vis_r4_o[6]));
assign Flf2z4 = (Jnf2z4 & Qnf2z4);
assign Qnf2z4 = (Xnf2z4 & Eof2z4);
assign Eof2z4 = (~(Fnd2z4 & vis_r1_o[6]));
assign Xnf2z4 = (~(Mnd2z4 & vis_r0_o[6]));
assign Jnf2z4 = (Lof2z4 & Sof2z4);
assign Sof2z4 = (~(Hod2z4 & vis_r3_o[6]));
assign Lof2z4 = (~(Ood2z4 & vis_r7_o[6]));
assign Jgf2z4 = (Zof2z4 & Gpf2z4);
assign Gpf2z4 = (~(Lpqvx4 & Zvqwx4));
assign Zvqwx4 = (!Bywwx4);
assign Bywwx4 = (Npf2z4 & Upf2z4);
assign Upf2z4 = (Bqf2z4 & Iqf2z4);
assign Iqf2z4 = (Pqf2z4 & Wqf2z4);
assign Wqf2z4 = (~(Nkd2z4 & vis_r2_o[7]));
assign Pqf2z4 = (~(Ukd2z4 & vis_r6_o[7]));
assign Bqf2z4 = (Drf2z4 & Krf2z4);
assign Krf2z4 = (~(Pld2z4 & vis_r5_o[7]));
assign Drf2z4 = (~(Wld2z4 & vis_r4_o[7]));
assign Npf2z4 = (Rrf2z4 & Yrf2z4);
assign Yrf2z4 = (Fsf2z4 & Msf2z4);
assign Msf2z4 = (~(Fnd2z4 & vis_r1_o[7]));
assign Fsf2z4 = (~(Mnd2z4 & vis_r0_o[7]));
assign Rrf2z4 = (Tsf2z4 & Atf2z4);
assign Atf2z4 = (~(Hod2z4 & vis_r3_o[7]));
assign Tsf2z4 = (~(Ood2z4 & vis_r7_o[7]));
assign Zof2z4 = (~(Onwwx4 & Xuqwx4));
assign Xuqwx4 = (!Lr9wx4);
assign Lr9wx4 = (Htf2z4 & Otf2z4);
assign Otf2z4 = (Vtf2z4 & Cuf2z4);
assign Cuf2z4 = (Juf2z4 & Quf2z4);
assign Quf2z4 = (~(Nkd2z4 & vis_r2_o[8]));
assign Juf2z4 = (~(Ukd2z4 & vis_r6_o[8]));
assign Vtf2z4 = (Xuf2z4 & Evf2z4);
assign Evf2z4 = (~(Pld2z4 & vis_r5_o[8]));
assign Xuf2z4 = (~(Wld2z4 & vis_r4_o[8]));
assign Htf2z4 = (Lvf2z4 & Svf2z4);
assign Svf2z4 = (Zvf2z4 & Gwf2z4);
assign Gwf2z4 = (~(Fnd2z4 & vis_r1_o[8]));
assign Zvf2z4 = (~(Mnd2z4 & vis_r0_o[8]));
assign Lvf2z4 = (Nwf2z4 & Uwf2z4);
assign Uwf2z4 = (~(Hod2z4 & vis_r3_o[8]));
assign Nwf2z4 = (~(Ood2z4 & vis_r7_o[8]));
assign Vff2z4 = (Bxf2z4 & Ixf2z4);
assign Ixf2z4 = (Pxf2z4 & Wxf2z4);
assign Wxf2z4 = (~(H9xvx4 & Ubqwx4));
assign Ubqwx4 = (!Duuwx4);
assign Duuwx4 = (Dyf2z4 & Kyf2z4);
assign Kyf2z4 = (Ryf2z4 & Yyf2z4);
assign Yyf2z4 = (Fzf2z4 & Mzf2z4);
assign Mzf2z4 = (~(vis_r2_o[1] & Nkd2z4));
assign Fzf2z4 = (~(vis_r6_o[1] & Ukd2z4));
assign Ryf2z4 = (Tzf2z4 & A0g2z4);
assign A0g2z4 = (~(vis_r5_o[1] & Pld2z4));
assign Tzf2z4 = (~(vis_r4_o[1] & Wld2z4));
assign Dyf2z4 = (H0g2z4 & O0g2z4);
assign O0g2z4 = (V0g2z4 & C1g2z4);
assign C1g2z4 = (~(vis_r1_o[1] & Fnd2z4));
assign V0g2z4 = (~(vis_r0_o[1] & Mnd2z4));
assign H0g2z4 = (J1g2z4 & Q1g2z4);
assign Q1g2z4 = (~(vis_r3_o[1] & Hod2z4));
assign J1g2z4 = (~(vis_r7_o[1] & Ood2z4));
assign Pxf2z4 = (~(Spqvx4 & Ituwx4));
assign Ituwx4 = (!Ylbwx4);
assign Ylbwx4 = (X1g2z4 & E2g2z4);
assign E2g2z4 = (L2g2z4 & S2g2z4);
assign S2g2z4 = (Z2g2z4 & G3g2z4);
assign G3g2z4 = (~(vis_r2_o[2] & Nkd2z4));
assign Z2g2z4 = (~(vis_r6_o[2] & Ukd2z4));
assign L2g2z4 = (N3g2z4 & U3g2z4);
assign U3g2z4 = (~(vis_r5_o[2] & Pld2z4));
assign N3g2z4 = (~(vis_r4_o[2] & Wld2z4));
assign X1g2z4 = (B4g2z4 & I4g2z4);
assign I4g2z4 = (P4g2z4 & W4g2z4);
assign W4g2z4 = (~(vis_r1_o[2] & Fnd2z4));
assign P4g2z4 = (~(vis_r0_o[2] & Mnd2z4));
assign B4g2z4 = (D5g2z4 & K5g2z4);
assign K5g2z4 = (~(vis_r3_o[2] & Hod2z4));
assign D5g2z4 = (~(vis_r7_o[2] & Ood2z4));
assign Bxf2z4 = (R5g2z4 & Y5g2z4);
assign Y5g2z4 = (~(Lpqvx4 & Iqqwx4));
assign Iqqwx4 = (!Ebbwx4);
assign Ebbwx4 = (F6g2z4 & M6g2z4);
assign M6g2z4 = (T6g2z4 & A7g2z4);
assign A7g2z4 = (H7g2z4 & O7g2z4);
assign O7g2z4 = (~(vis_r2_o[3] & Nkd2z4));
assign H7g2z4 = (~(vis_r6_o[3] & Ukd2z4));
assign T6g2z4 = (V7g2z4 & C8g2z4);
assign C8g2z4 = (~(vis_r5_o[3] & Pld2z4));
assign V7g2z4 = (~(vis_r4_o[3] & Wld2z4));
assign F6g2z4 = (J8g2z4 & Q8g2z4);
assign Q8g2z4 = (X8g2z4 & E9g2z4);
assign E9g2z4 = (~(vis_r1_o[3] & Fnd2z4));
assign X8g2z4 = (~(vis_r0_o[3] & Mnd2z4));
assign J8g2z4 = (L9g2z4 & S9g2z4);
assign S9g2z4 = (~(vis_r3_o[3] & Hod2z4));
assign L9g2z4 = (~(vis_r7_o[3] & Ood2z4));
assign R5g2z4 = (~(Onwwx4 & Drqwx4));
assign Drqwx4 = (!Bdwwx4);
assign Bdwwx4 = (Z9g2z4 & Gag2z4);
assign Gag2z4 = (Nag2z4 & Uag2z4);
assign Uag2z4 = (Bbg2z4 & Ibg2z4);
assign Ibg2z4 = (~(vis_r2_o[4] & Nkd2z4));
assign Bbg2z4 = (~(vis_r6_o[4] & Ukd2z4));
assign Nag2z4 = (Pbg2z4 & Wbg2z4);
assign Wbg2z4 = (~(vis_r5_o[4] & Pld2z4));
assign Pbg2z4 = (~(vis_r4_o[4] & Wld2z4));
assign Z9g2z4 = (Dcg2z4 & Kcg2z4);
assign Kcg2z4 = (Rcg2z4 & Ycg2z4);
assign Ycg2z4 = (~(vis_r1_o[4] & Fnd2z4));
assign Rcg2z4 = (~(vis_r0_o[4] & Mnd2z4));
assign Dcg2z4 = (Fdg2z4 & Mdg2z4);
assign Mdg2z4 = (~(vis_r3_o[4] & Hod2z4));
assign Fdg2z4 = (~(vis_r7_o[4] & Ood2z4));
assign Hff2z4 = (Yryvx4 ? Aeg2z4 : Tdg2z4);
assign Yryvx4 = (!Qm9vx4);
assign Aeg2z4 = (Heg2z4 & Oeg2z4);
assign Oeg2z4 = (Veg2z4 & Cfg2z4);
assign Cfg2z4 = (~(H9xvx4 & Niqwx4));
assign Niqwx4 = (!Zkuwx4);
assign Zkuwx4 = (Jfg2z4 & Qfg2z4);
assign Qfg2z4 = (Xfg2z4 & Egg2z4);
assign Egg2z4 = (Lgg2z4 & Sgg2z4);
assign Sgg2z4 = (~(Nkd2z4 & vis_r2_o[13]));
assign Lgg2z4 = (~(Ukd2z4 & vis_r6_o[13]));
assign Xfg2z4 = (Zgg2z4 & Ghg2z4);
assign Ghg2z4 = (~(Pld2z4 & vis_r5_o[13]));
assign Zgg2z4 = (~(Wld2z4 & vis_r4_o[13]));
assign Jfg2z4 = (Nhg2z4 & Uhg2z4);
assign Uhg2z4 = (Big2z4 & Iig2z4);
assign Iig2z4 = (~(Fnd2z4 & vis_r1_o[13]));
assign Big2z4 = (~(Mnd2z4 & vis_r0_o[13]));
assign Nhg2z4 = (Pig2z4 & Wig2z4);
assign Wig2z4 = (~(Hod2z4 & vis_r3_o[13]));
assign Pig2z4 = (~(Ood2z4 & vis_r7_o[13]));
assign Veg2z4 = (~(Spqvx4 & Uluwx4));
assign Uluwx4 = (!Hmqwx4);
assign Hmqwx4 = (Djg2z4 & Kjg2z4);
assign Kjg2z4 = (Rjg2z4 & Yjg2z4);
assign Yjg2z4 = (Fkg2z4 & Mkg2z4);
assign Mkg2z4 = (~(Nkd2z4 & vis_r2_o[14]));
assign Fkg2z4 = (~(Ukd2z4 & vis_r6_o[14]));
assign Rjg2z4 = (Tkg2z4 & Alg2z4);
assign Alg2z4 = (~(Pld2z4 & vis_r5_o[14]));
assign Tkg2z4 = (~(Wld2z4 & vis_r4_o[14]));
assign Djg2z4 = (Hlg2z4 & Olg2z4);
assign Olg2z4 = (Vlg2z4 & Cmg2z4);
assign Cmg2z4 = (~(Fnd2z4 & vis_r1_o[14]));
assign Vlg2z4 = (~(Mnd2z4 & vis_r0_o[14]));
assign Hlg2z4 = (Jmg2z4 & Qmg2z4);
assign Qmg2z4 = (~(Hod2z4 & vis_r3_o[14]));
assign Jmg2z4 = (~(Ood2z4 & vis_r7_o[14]));
assign Heg2z4 = (Xmg2z4 & Eng2z4);
assign Eng2z4 = (~(Lpqvx4 & Omqwx4));
assign Omqwx4 = (!Ey9wx4);
assign Ey9wx4 = (Lng2z4 & Sng2z4);
assign Sng2z4 = (Zng2z4 & Gog2z4);
assign Gog2z4 = (Nog2z4 & Uog2z4);
assign Uog2z4 = (~(Nkd2z4 & vis_r2_o[15]));
assign Nog2z4 = (~(Ukd2z4 & vis_r6_o[15]));
assign Zng2z4 = (Bpg2z4 & Ipg2z4);
assign Ipg2z4 = (~(Pld2z4 & vis_r5_o[15]));
assign Bpg2z4 = (~(Wld2z4 & vis_r4_o[15]));
assign Lng2z4 = (Ppg2z4 & Wpg2z4);
assign Wpg2z4 = (Dqg2z4 & Kqg2z4);
assign Kqg2z4 = (~(Fnd2z4 & vis_r1_o[15]));
assign Dqg2z4 = (~(Mnd2z4 & vis_r0_o[15]));
assign Ppg2z4 = (Rqg2z4 & Yqg2z4);
assign Yqg2z4 = (~(Hod2z4 & vis_r3_o[15]));
assign Rqg2z4 = (~(Ood2z4 & vis_r7_o[15]));
assign Xmg2z4 = (~(Onwwx4 & Mlqwx4));
assign Mlqwx4 = (!Nrvwx4);
assign Nrvwx4 = (Frg2z4 & Mrg2z4);
assign Mrg2z4 = (Trg2z4 & Asg2z4);
assign Asg2z4 = (Hsg2z4 & Osg2z4);
assign Osg2z4 = (~(Nkd2z4 & vis_r2_o[16]));
assign Hsg2z4 = (~(Ukd2z4 & vis_r6_o[16]));
assign Trg2z4 = (Vsg2z4 & Ctg2z4);
assign Ctg2z4 = (~(Pld2z4 & vis_r5_o[16]));
assign Vsg2z4 = (~(Wld2z4 & vis_r4_o[16]));
assign Frg2z4 = (Jtg2z4 & Qtg2z4);
assign Qtg2z4 = (Xtg2z4 & Eug2z4);
assign Eug2z4 = (~(Fnd2z4 & vis_r1_o[16]));
assign Xtg2z4 = (~(Mnd2z4 & vis_r0_o[16]));
assign Jtg2z4 = (Lug2z4 & Sug2z4);
assign Sug2z4 = (~(Hod2z4 & vis_r3_o[16]));
assign Lug2z4 = (~(Ood2z4 & vis_r7_o[16]));
assign Tdg2z4 = (Zug2z4 & Gvg2z4);
assign Gvg2z4 = (Nvg2z4 & Uvg2z4);
assign Uvg2z4 = (~(H9xvx4 & Quqwx4));
assign Quqwx4 = (!Pybwx4);
assign Pybwx4 = (Bwg2z4 & Iwg2z4);
assign Iwg2z4 = (Pwg2z4 & Wwg2z4);
assign Wwg2z4 = (Dxg2z4 & Kxg2z4);
assign Kxg2z4 = (~(vis_r2_o[9] & Nkd2z4));
assign Dxg2z4 = (~(vis_r6_o[9] & Ukd2z4));
assign Pwg2z4 = (Rxg2z4 & Yxg2z4);
assign Yxg2z4 = (~(vis_r5_o[9] & Pld2z4));
assign Rxg2z4 = (~(vis_r4_o[9] & Wld2z4));
assign Bwg2z4 = (Fyg2z4 & Myg2z4);
assign Myg2z4 = (Tyg2z4 & Azg2z4);
assign Azg2z4 = (~(vis_r1_o[9] & Fnd2z4));
assign Tyg2z4 = (~(vis_r0_o[9] & Mnd2z4));
assign Fyg2z4 = (Hzg2z4 & Ozg2z4);
assign Ozg2z4 = (~(vis_r3_o[9] & Hod2z4));
assign Hzg2z4 = (~(vis_r7_o[9] & Ood2z4));
assign H9xvx4 = (Ik9vx4 & Ml9vx4);
assign Nvg2z4 = (~(Spqvx4 & I0vwx4));
assign I0vwx4 = (!Pjqwx4);
assign Pjqwx4 = (Vzg2z4 & C0h2z4);
assign C0h2z4 = (J0h2z4 & Q0h2z4);
assign Q0h2z4 = (X0h2z4 & E1h2z4);
assign E1h2z4 = (~(vis_r2_o[10] & Nkd2z4));
assign X0h2z4 = (~(vis_r6_o[10] & Ukd2z4));
assign J0h2z4 = (L1h2z4 & S1h2z4);
assign S1h2z4 = (~(vis_r5_o[10] & Pld2z4));
assign L1h2z4 = (~(vis_r4_o[10] & Wld2z4));
assign Vzg2z4 = (Z1h2z4 & G2h2z4);
assign G2h2z4 = (N2h2z4 & U2h2z4);
assign U2h2z4 = (~(vis_r1_o[10] & Fnd2z4));
assign N2h2z4 = (~(vis_r0_o[10] & Mnd2z4));
assign Z1h2z4 = (B3h2z4 & I3h2z4);
assign I3h2z4 = (~(vis_r3_o[10] & Hod2z4));
assign B3h2z4 = (~(vis_r7_o[10] & Ood2z4));
assign Spqvx4 = (~(P3h2z4 | Ik9vx4));
assign Zug2z4 = (W3h2z4 & D4h2z4);
assign D4h2z4 = (~(Lpqvx4 & Uiqwx4));
assign Uiqwx4 = (!Ai9wx4);
assign Ai9wx4 = (K4h2z4 & R4h2z4);
assign R4h2z4 = (Y4h2z4 & F5h2z4);
assign F5h2z4 = (M5h2z4 & T5h2z4);
assign T5h2z4 = (~(Nkd2z4 & vis_r2_o[11]));
assign M5h2z4 = (~(Ukd2z4 & vis_r6_o[11]));
assign Y4h2z4 = (A6h2z4 & H6h2z4);
assign H6h2z4 = (~(Pld2z4 & vis_r5_o[11]));
assign A6h2z4 = (~(Wld2z4 & vis_r4_o[11]));
assign K4h2z4 = (O6h2z4 & V6h2z4);
assign V6h2z4 = (C7h2z4 & J7h2z4);
assign J7h2z4 = (~(Fnd2z4 & vis_r1_o[11]));
assign C7h2z4 = (~(Mnd2z4 & vis_r0_o[11]));
assign O6h2z4 = (Q7h2z4 & X7h2z4);
assign X7h2z4 = (~(Hod2z4 & vis_r3_o[11]));
assign Q7h2z4 = (~(Ood2z4 & vis_r7_o[11]));
assign Lpqvx4 = (~(Cppvx4 | Ml9vx4));
assign W3h2z4 = (~(Onwwx4 & Wjqwx4));
assign Wjqwx4 = (!H2wwx4);
assign H2wwx4 = (E8h2z4 & L8h2z4);
assign L8h2z4 = (S8h2z4 & Z8h2z4);
assign Z8h2z4 = (G9h2z4 & N9h2z4);
assign N9h2z4 = (~(Nkd2z4 & vis_r2_o[12]));
assign Nkd2z4 = (~(U9h2z4 | Erc2z4));
assign G9h2z4 = (~(Ukd2z4 & vis_r6_o[12]));
assign Ukd2z4 = (~(Bah2z4 | Erc2z4));
assign Erc2z4 = (~(Tjh2z4[1] & Iah2z4));
assign S8h2z4 = (Pah2z4 & Wah2z4);
assign Wah2z4 = (~(Pld2z4 & vis_r5_o[12]));
assign Pld2z4 = (~(Ptc2z4 | Bah2z4));
assign Pah2z4 = (~(Wld2z4 & vis_r4_o[12]));
assign Wld2z4 = (~(Lrc2z4 | Bah2z4));
assign E8h2z4 = (Dbh2z4 & Kbh2z4);
assign Kbh2z4 = (Rbh2z4 & Ybh2z4);
assign Ybh2z4 = (~(Fnd2z4 & vis_r1_o[12]));
assign Fnd2z4 = (~(Ptc2z4 | U9h2z4));
assign Ptc2z4 = (!Mja2z4);
assign Mja2z4 = (Tjh2z4[0] & Fch2z4);
assign Rbh2z4 = (~(Mnd2z4 & vis_r0_o[12]));
assign Mnd2z4 = (~(Lrc2z4 | U9h2z4));
assign Lrc2z4 = (~(Iah2z4 & Fch2z4));
assign Fch2z4 = (!Tjh2z4[1]);
assign Iah2z4 = (!Tjh2z4[0]);
assign Dbh2z4 = (Mch2z4 & Tch2z4);
assign Tch2z4 = (~(Hod2z4 & vis_r3_o[12]));
assign Hod2z4 = (~(U9h2z4 | Nsc2z4));
assign U9h2z4 = (Tjh2z4[2] | Tjh2z4[3]);
assign Mch2z4 = (~(Ood2z4 & vis_r7_o[12]));
assign Ood2z4 = (~(Bah2z4 | Nsc2z4));
assign Nsc2z4 = (~(Tjh2z4[1] & Tjh2z4[0]));
assign Bah2z4 = (~(Tjh2z4[2] & Wtc2z4));
assign Wtc2z4 = (!Tjh2z4[3]);
assign Onwwx4 = (Cppvx4 & P3h2z4);
assign P3h2z4 = (!Ml9vx4);
assign Cppvx4 = (!Ik9vx4);
assign Wed2z4 = (S87wx4 | W5yvx4);
assign S87wx4 = (!Ncqvx4);
assign Ncqvx4 = (~(Us2wx4 | Mcgvx4));
assign Ied2z4 = (Whgvx4 & Adh2z4);
assign Adh2z4 = (M93wx4 | B1ovx4);
assign M93wx4 = (!X77wx4);
assign X77wx4 = (Mcgvx4 & U9gvx4);
assign Oq42z4 = (Qr42z4 & Hdh2z4);
assign Hdh2z4 = (~(Odh2z4 & Vdh2z4));
assign Vdh2z4 = (Fpfwx4 | Efgvx4);
assign Fpfwx4 = (!Kngwx4);
assign Kngwx4 = (Nggvx4 & F3ovx4);
assign Odh2z4 = (~(R5dwx4 | H5mwx4));
assign H5mwx4 = (~(F3ovx4 | Us2wx4));
assign F3ovx4 = (!Z6gvx4);
assign R5dwx4 = (~(U9gvx4 | Efgvx4));
assign Qr42z4 = (Ceh2z4 & Jeh2z4);
assign Jeh2z4 = (Qeh2z4 & Z2dwx4);
assign Z2dwx4 = (!Liiwx4);
assign Liiwx4 = (~(U9gvx4 | Dbgvx4));
assign Qeh2z4 = (~(Xeh2z4 & Nggvx4));
assign Xeh2z4 = (U9gvx4 & Hw2wx4);
assign Hw2wx4 = (~(Us2wx4 | B1ovx4));
assign B1ovx4 = (!Dbgvx4);
assign Us2wx4 = (!Efgvx4);
assign Ceh2z4 = (Efh2z4 & Lfh2z4);
assign Lfh2z4 = (E78wx4 | T93wx4);
assign T93wx4 = (!Socwx4);
assign Socwx4 = (~(U0ovx4 | Efgvx4));
assign U0ovx4 = (!Whgvx4);
assign E78wx4 = (!Fhc2z4);
assign Fhc2z4 = (~(W5yvx4 | U9gvx4));
assign W5yvx4 = (!Nggvx4);
assign Efh2z4 = (Mcgvx4 | Cn8vx4);

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J6i2z4 <= 1'b0;
  else
    J6i2z4 <= Elnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z7i2z4 <= 1'b1;
  else
    Z7i2z4 <= Ojnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H9i2z4 <= 1'b1;
  else
    H9i2z4 <= M4nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wai2z4 <= 1'b1;
  else
    Wai2z4 <= Lyhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gci2z4 <= 1'b1;
  else
    Gci2z4 <= V3ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pdi2z4 <= 1'b1;
  else
    Pdi2z4 <= Eyhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zei2z4 <= 1'b0;
  else
    Zei2z4 <= Finvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Igi2z4 <= 1'b1;
  else
    Igi2z4 <= Cflvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rhi2z4 <= 1'b1;
  else
    Rhi2z4 <= Velvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gji2z4 <= 1'b0;
  else
    Gji2z4 <= H3ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tki2z4 <= 1'b0;
  else
    Tki2z4 <= Xxhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Emi2z4 <= 1'b0;
  else
    Emi2z4 <= Qxhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rni2z4 <= 1'b1;
  else
    Rni2z4 <= Jxhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fpi2z4 <= 1'b1;
  else
    Fpi2z4 <= B7ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uqi2z4 <= 1'b0;
  else
    Uqi2z4 <= Mcmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Isi2z4 <= 1'b1;
  else
    Isi2z4 <= Frlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xti2z4 <= 1'b1;
  else
    Xti2z4 <= Wgnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mvi2z4 <= 1'b0;
  else
    Mvi2z4 <= E8mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ywi2z4 <= 1'b0;
  else
    Ywi2z4 <= Owgvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kyi2z4 <= 1'b1;
  else
    Kyi2z4 <= Vcnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yzi2z4 <= 1'b1;
  else
    Yzi2z4 <= Qdnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M1j2z4 <= 1'b1;
  else
    M1j2z4 <= Hllvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X2j2z4 <= 1'b1;
  else
    X2j2z4 <= Rjlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M4j2z4 <= 1'b1;
  else
    M4j2z4 <= W7ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B6j2z4 <= 1'b1;
  else
    B6j2z4 <= K8ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q7j2z4 <= 1'b1;
  else
    Q7j2z4 <= Vjnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F9j2z4 <= 1'b1;
  else
    F9j2z4 <= Lvkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uaj2z4 <= 1'b0;
  else
    Uaj2z4 <= U9mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fcj2z4 <= 1'b1;
  else
    Fcj2z4 <= Cxhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qdj2z4 <= 1'b1;
  else
    Qdj2z4 <= Llnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ffj2z4 <= 1'b0;
  else
    Ffj2z4 <= Vwhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sgj2z4 <= 1'b0;
  else
    Sgj2z4 <= Owhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fij2z4 <= 1'b0;
  else
    Fij2z4 <= Hwhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sjj2z4 <= 1'b1;
  else
    Sjj2z4 <= Awhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Glj2z4 <= 1'b1;
  else
    Glj2z4 <= Nolvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vmj2z4 <= 1'b1;
  else
    Vmj2z4 <= Xukvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Koj2z4 <= 1'b1;
  else
    Koj2z4 <= Gfnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zpj2z4 <= 1'b1;
  else
    Zpj2z4 <= Tskvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Orj2z4 <= 1'b1;
  else
    Orj2z4 <= J4ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dtj2z4 <= 1'b1;
  else
    Dtj2z4 <= Snlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ruj2z4 <= 1'b1;
  else
    Ruj2z4 <= Kqlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fwj2z4 <= 1'b1;
  else
    Fwj2z4 <= Lenvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Txj2z4 <= 1'b1;
  else
    Txj2z4 <= Minvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hzj2z4 <= 1'b0;
  else
    Hzj2z4 <= M5mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V0k2z4 <= 1'b1;
  else
    V0k2z4 <= Q1lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K2k2z4 <= 1'b1;
  else
    K2k2z4 <= U3lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z3k2z4 <= 1'b1;
  else
    Z3k2z4 <= I4lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O5k2z4 <= 1'b1;
  else
    O5k2z4 <= D5lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D7k2z4 <= 1'b1;
  else
    D7k2z4 <= K5lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S8k2z4 <= 1'b1;
  else
    S8k2z4 <= R5lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hak2z4 <= 1'b1;
  else
    Hak2z4 <= Galvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wbk2z4 <= 1'b0;
  else
    Wbk2z4 <= T5mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Idk2z4 <= 1'b0;
  else
    Idk2z4 <= Rhnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rek2z4 <= 1'b1;
  else
    Rek2z4 <= Yjlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ggk2z4 <= 1'b1;
  else
    Ggk2z4 <= Golvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vhk2z4 <= 1'b1;
  else
    Vhk2z4 <= Yqlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kjk2z4 <= 1'b1;
  else
    Kjk2z4 <= Zenvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zkk2z4 <= 1'b1;
  else
    Zkk2z4 <= Dhnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Omk2z4 <= 1'b1;
  else
    Omk2z4 <= Tvhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aok2z4 <= 1'b0;
  else
    Aok2z4 <= Mvhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Npk2z4 <= 1'b0;
  else
    Npk2z4 <= Fvhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ark2z4 <= 1'b0;
  else
    Ark2z4 <= Yuhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nsk2z4 <= 1'b0;
  else
    Nsk2z4 <= Ruhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Auk2z4 <= 1'b1;
  else
    Auk2z4 <= P3mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Svk2z4 <= 1'b1;
  else
    Svk2z4 <= Kuhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gxk2z4 <= 1'b0;
  else
    Gxk2z4 <= T2ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xyk2z4 <= 1'b1;
  else
    Xyk2z4 <= Duhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J0l2z4 <= 1'b1;
  else
    J0l2z4 <= Wthvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V1l2z4 <= 1'b1;
  else
    V1l2z4 <= O3ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K3l2z4 <= 1'b0;
  else
    K3l2z4 <= F4nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z4l2z4 <= 1'b0;
  else
    Z4l2z4 <= Bhmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q6l2z4 <= 1'b0;
  else
    Q6l2z4 <= Ugmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H8l2z4 <= 1'b0;
  else
    H8l2z4 <= Ngmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y9l2z4 <= 1'b0;
  else
    Y9l2z4 <= I0ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pbl2z4 <= 1'b1;
  else
    Pbl2z4 <= Bxkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Edl2z4 <= 1'b1;
  else
    Edl2z4 <= Fzkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tel2z4 <= 1'b1;
  else
    Tel2z4 <= Tzkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Igl2z4 <= 1'b1;
  else
    Igl2z4 <= O0lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xhl2z4 <= 1'b1;
  else
    Xhl2z4 <= V0lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mjl2z4 <= 1'b0;
  else
    Mjl2z4 <= Nmnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cll2z4 <= 1'b1;
  else
    Cll2z4 <= Fklvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qml2z4 <= 1'b1;
  else
    Qml2z4 <= Znlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eol2z4 <= 1'b1;
  else
    Eol2z4 <= Rqlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Spl2z4 <= 1'b1;
  else
    Spl2z4 <= Senvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Grl2z4 <= 1'b1;
  else
    Grl2z4 <= Ignvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Usl2z4 <= 1'b0;
  else
    Usl2z4 <= Phmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lul2z4 <= 1'b0;
  else
    Lul2z4 <= Syhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dwl2z4 <= 1'b1;
  else
    Dwl2z4 <= Hcnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rxl2z4 <= 1'b1;
  else
    Rxl2z4 <= S7nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fzl2z4 <= 1'b1;
  else
    Fzl2z4 <= Jdnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T0m2z4 <= 1'b1;
  else
    T0m2z4 <= Lakvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H2m2z4 <= 1'b1;
  else
    H2m2z4 <= Pckvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V3m2z4 <= 1'b1;
  else
    V3m2z4 <= Ddkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J5m2z4 <= 1'b1;
  else
    J5m2z4 <= Ydkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X6m2z4 <= 1'b1;
  else
    X6m2z4 <= Fekvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L8m2z4 <= 1'b1;
  else
    L8m2z4 <= Gumvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cam2z4 <= 1'b0;
  else
    Cam2z4 <= L8mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nbm2z4 <= 1'b0;
  else
    Nbm2z4 <= Zlnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bdm2z4 <= 1'b1;
  else
    Bdm2z4 <= U8nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qem2z4 <= 1'b1;
  else
    Qem2z4 <= Ajnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fgm2z4 <= 1'b1;
  else
    Fgm2z4 <= Pthvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Thm2z4 <= 1'b0;
  else
    Thm2z4 <= Xdnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ejm2z4 <= 1'b1;
  else
    Ejm2z4 <= Lnlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Skm2z4 <= 1'b1;
  else
    Skm2z4 <= Dqlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gmm2z4 <= 1'b1;
  else
    Gmm2z4 <= Eenvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Unm2z4 <= 1'b1;
  else
    Unm2z4 <= Bgnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ipm2z4 <= 1'b1;
  else
    Ipm2z4 <= Eokvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wqm2z4 <= 1'b1;
  else
    Wqm2z4 <= Iqkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ksm2z4 <= 1'b1;
  else
    Ksm2z4 <= Wqkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ytm2z4 <= 1'b1;
  else
    Ytm2z4 <= Rrkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mvm2z4 <= 1'b1;
  else
    Mvm2z4 <= Yrkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Axm2z4 <= 1'b0;
  else
    Axm2z4 <= Whmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rym2z4 <= 1'b0;
  else
    Rym2z4 <= Zyhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J0n2z4 <= 1'b1;
  else
    J0n2z4 <= P5kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y1n2z4 <= 1'b1;
  else
    Y1n2z4 <= T7kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N3n2z4 <= 1'b1;
  else
    N3n2z4 <= H8kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C5n2z4 <= 1'b1;
  else
    C5n2z4 <= C9kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R6n2z4 <= 1'b1;
  else
    R6n2z4 <= J9kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G8n2z4 <= 1'b0;
  else
    G8n2z4 <= Ihmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X9n2z4 <= 1'b0;
  else
    X9n2z4 <= Tcmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lbn2z4 <= 1'b1;
  else
    Lbn2z4 <= Tbnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zcn2z4 <= 1'b1;
  else
    Zcn2z4 <= U2mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nen2z4 <= 1'b0;
  else
    Nen2z4 <= Ollvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yfn2z4 <= 1'b1;
  else
    Yfn2z4 <= Rmivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mhn2z4 <= 1'b1;
  else
    Mhn2z4 <= Voivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ajn2z4 <= 1'b1;
  else
    Ajn2z4 <= Jpivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Okn2z4 <= 1'b1;
  else
    Okn2z4 <= Eqivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cmn2z4 <= 1'b1;
  else
    Cmn2z4 <= Lqivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qnn2z4 <= 1'b0;
  else
    Qnn2z4 <= C7mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ipn2z4 <= 1'b0;
  else
    Ipn2z4 <= B0ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Arn2z4 <= 1'b1;
  else
    Arn2z4 <= Hnjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Psn2z4 <= 1'b1;
  else
    Psn2z4 <= Lpjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eun2z4 <= 1'b1;
  else
    Eun2z4 <= Zpjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tvn2z4 <= 1'b1;
  else
    Tvn2z4 <= Uqjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ixn2z4 <= 1'b1;
  else
    Ixn2z4 <= Brjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xyn2z4 <= 1'b1;
  else
    Xyn2z4 <= Numvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O0o2z4 <= 1'b1;
  else
    O0o2z4 <= Iomvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F2o2z4 <= 1'b1;
  else
    F2o2z4 <= Etmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V3o2z4 <= 1'b0;
  else
    V3o2z4 <= Rbmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J5o2z4 <= 1'b1;
  else
    J5o2z4 <= Dejvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y6o2z4 <= 1'b1;
  else
    Y6o2z4 <= Hgjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N8o2z4 <= 1'b1;
  else
    N8o2z4 <= Vgjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cao2z4 <= 1'b1;
  else
    Cao2z4 <= Qhjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rbo2z4 <= 1'b1;
  else
    Rbo2z4 <= Xhjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gdo2z4 <= 1'b1;
  else
    Gdo2z4 <= Bvmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xeo2z4 <= 1'b1;
  else
    Xeo2z4 <= Womvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ogo2z4 <= 1'b1;
  else
    Ogo2z4 <= Nnmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fio2z4 <= 1'b1;
  else
    Fio2z4 <= Ualvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ujo2z4 <= 1'b1;
  else
    Ujo2z4 <= Yclvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jlo2z4 <= 1'b1;
  else
    Jlo2z4 <= Mdlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ymo2z4 <= 1'b1;
  else
    Ymo2z4 <= Helvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Noo2z4 <= 1'b1;
  else
    Noo2z4 <= Oelvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cqo2z4 <= 1'b1;
  else
    Cqo2z4 <= Yhnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rro2z4 <= 1'b1;
  else
    Rro2z4 <= Qflvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gto2z4 <= 1'b1;
  else
    Gto2z4 <= Uhlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vuo2z4 <= 1'b1;
  else
    Vuo2z4 <= Iilvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kwo2z4 <= 1'b1;
  else
    Kwo2z4 <= Sijvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zxo2z4 <= 1'b1;
  else
    Zxo2z4 <= Wkjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ozo2z4 <= 1'b1;
  else
    Ozo2z4 <= Kljvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D1p2z4 <= 1'b1;
  else
    D1p2z4 <= Fmjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S2p2z4 <= 1'b1;
  else
    S2p2z4 <= Mmjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H4p2z4 <= 1'b1;
  else
    H4p2z4 <= Tmjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W5p2z4 <= 1'b1;
  else
    W5p2z4 <= Irjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L7p2z4 <= 1'b1;
  else
    L7p2z4 <= Xvjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A9p2z4 <= 1'b1;
  else
    A9p2z4 <= Wrjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pap2z4 <= 1'b1;
  else
    Pap2z4 <= Aujvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ecp2z4 <= 1'b1;
  else
    Ecp2z4 <= Oujvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tdp2z4 <= 1'b0;
  else
    Tdp2z4 <= Wamvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Efp2z4 <= 1'b1;
  else
    Efp2z4 <= Qnkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sgp2z4 <= 1'b1;
  else
    Sgp2z4 <= Pjkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gip2z4 <= 1'b1;
  else
    Gip2z4 <= Tlkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ujp2z4 <= 1'b1;
  else
    Ujp2z4 <= Hmkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ilp2z4 <= 1'b1;
  else
    Ilp2z4 <= Cnkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wmp2z4 <= 1'b1;
  else
    Wmp2z4 <= Jnkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kop2z4 <= 1'b0;
  else
    Kop2z4 <= Xknvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aqp2z4 <= 1'b0;
  else
    Aqp2z4 <= Fcmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qrp2z4 <= 1'b0;
  else
    Qrp2z4 <= Ybmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gtp2z4 <= 1'b1;
  else
    Gtp2z4 <= Mbnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uup2z4 <= 1'b1;
  else
    Uup2z4 <= N2mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Iwp2z4 <= 1'b1;
  else
    Iwp2z4 <= D4mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wxp2z4 <= 1'b0;
  else
    Wxp2z4 <= X9kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mzp2z4 <= 1'b1;
  else
    Mzp2z4 <= O9jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B1q2z4 <= 1'b1;
  else
    B1q2z4 <= Sbjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q2q2z4 <= 1'b1;
  else
    Q2q2z4 <= Gcjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F4q2z4 <= 1'b1;
  else
    F4q2z4 <= Bdjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U5q2z4 <= 1'b1;
  else
    U5q2z4 <= Idjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J7q2z4 <= 1'b1;
  else
    J7q2z4 <= Pdjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y8q2z4 <= 1'b1;
  else
    Y8q2z4 <= Zcivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Naq2z4 <= 1'b1;
  else
    Naq2z4 <= Y8ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ccq2z4 <= 1'b1;
  else
    Ccq2z4 <= Cbivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rdq2z4 <= 1'b1;
  else
    Rdq2z4 <= Qbivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gfq2z4 <= 1'b1;
  else
    Gfq2z4 <= F6lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vgq2z4 <= 1'b1;
  else
    Vgq2z4 <= J8lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kiq2z4 <= 1'b1;
  else
    Kiq2z4 <= X8lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zjq2z4 <= 1'b1;
  else
    Zjq2z4 <= Ithvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Llq2z4 <= 1'b1;
  else
    Llq2z4 <= B5kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Anq2z4 <= 1'b1;
  else
    Anq2z4 <= A1kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Poq2z4 <= 1'b1;
  else
    Poq2z4 <= E3kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eqq2z4 <= 1'b1;
  else
    Eqq2z4 <= S3kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Trq2z4 <= 1'b0;
  else
    Trq2z4 <= Pamvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Etq2z4 <= 1'b0;
  else
    Etq2z4 <= Dbmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wuq2z4 <= 1'b0;
  else
    Wuq2z4 <= Gzhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Owq2z4 <= 1'b1;
  else
    Owq2z4 <= Fbnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cyq2z4 <= 1'b1;
  else
    Cyq2z4 <= Bthvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qzq2z4 <= 1'b1;
  else
    Qzq2z4 <= Tinvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E1r2z4 <= 1'b1;
  else
    E1r2z4 <= Afkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S2r2z4 <= 1'b1;
  else
    S2r2z4 <= Ehkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G4r2z4 <= 1'b1;
  else
    G4r2z4 <= Shkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U5r2z4 <= 1'b1;
  else
    U5r2z4 <= Nikvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I7r2z4 <= 1'b1;
  else
    I7r2z4 <= Uikvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W8r2z4 <= 1'b0;
  else
    W8r2z4 <= A6mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oar2z4 <= 1'b0;
  else
    Oar2z4 <= Nzhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gcr2z4 <= 1'b1;
  else
    Gcr2z4 <= K0jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vdr2z4 <= 1'b1;
  else
    Vdr2z4 <= O2jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kfr2z4 <= 1'b1;
  else
    Kfr2z4 <= C3jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zgr2z4 <= 1'b1;
  else
    Zgr2z4 <= X3jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oir2z4 <= 1'b1;
  else
    Oir2z4 <= E4jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dkr2z4 <= 1'b1;
  else
    Dkr2z4 <= L4jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Slr2z4 <= 1'b1;
  else
    Slr2z4 <= A9jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hnr2z4 <= 1'b1;
  else
    Hnr2z4 <= Z4jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wor2z4 <= 1'b1;
  else
    Wor2z4 <= D7jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lqr2z4 <= 1'b1;
  else
    Lqr2z4 <= R7jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Asr2z4 <= 1'b1;
  else
    Asr2z4 <= Ndivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Otr2z4 <= 1'b1;
  else
    Otr2z4 <= Rfivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cvr2z4 <= 1'b1;
  else
    Cvr2z4 <= Fgivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qwr2z4 <= 1'b1;
  else
    Qwr2z4 <= Ahivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eyr2z4 <= 1'b1;
  else
    Eyr2z4 <= Hhivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Szr2z4 <= 1'b1;
  else
    Szr2z4 <= Ohivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G1s2z4 <= 1'b1;
  else
    G1s2z4 <= Dmivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U2s2z4 <= 1'b1;
  else
    U2s2z4 <= Ciivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I4s2z4 <= 1'b1;
  else
    I4s2z4 <= Gkivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W5s2z4 <= 1'b1;
  else
    W5s2z4 <= Ukivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K7s2z4 <= 1'b1;
  else
    K7s2z4 <= Grivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z8s2z4 <= 1'b1;
  else
    Z8s2z4 <= Ktivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oas2z4 <= 1'b1;
  else
    Oas2z4 <= Ytivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dcs2z4 <= 1'b1;
  else
    Dcs2z4 <= Tuivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rds2z4 <= 1'b1;
  else
    Rds2z4 <= Avivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ffs2z4 <= 1'b0;
  else
    Ffs2z4 <= Qknvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vgs2z4 <= 1'b0;
  else
    Vgs2z4 <= Xlmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mis2z4 <= 1'b0;
  else
    Mis2z4 <= Emmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dks2z4 <= 1'b0;
  else
    Dks2z4 <= Qlmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uls2z4 <= 1'b0;
  else
    Uls2z4 <= Jlmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lns2z4 <= 1'b0;
  else
    Lns2z4 <= Clmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cps2z4 <= 1'b0;
  else
    Cps2z4 <= Vkmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tqs2z4 <= 1'b0;
  else
    Tqs2z4 <= Tjmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kss2z4 <= 1'b0;
  else
    Kss2z4 <= Akmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bus2z4 <= 1'b0;
  else
    Bus2z4 <= Mjmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Svs2z4 <= 1'b0;
  else
    Svs2z4 <= Fjmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jxs2z4 <= 1'b0;
  else
    Jxs2z4 <= Yimvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Azs2z4 <= 1'b0;
  else
    Azs2z4 <= Rimvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R0t2z4 <= 1'b0;
  else
    R0t2z4 <= Odmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I2t2z4 <= 1'b1;
  else
    I2t2z4 <= W3mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A4t2z4 <= 1'b0;
  else
    A4t2z4 <= Nfnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O5t2z4 <= 1'b1;
  else
    O5t2z4 <= Ushvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y6t2z4 <= 1'b0;
  else
    Y6t2z4 <= Nshvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L8t2z4 <= 1'b0;
  else
    L8t2z4 <= Cdnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y9t2z4 <= 1'b0;
  else
    Y9t2z4 <= Gshvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mbt2z4 <= 1'b0;
  else
    Mbt2z4 <= Vdmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Adt2z4 <= 1'b0;
  else
    Adt2z4 <= Cemvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pet2z4 <= 1'b0;
  else
    Pet2z4 <= Zrhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cgt2z4 <= 1'b1;
  else
    Cgt2z4 <= Wplvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rht2z4 <= 1'b1;
  else
    Rht2z4 <= Pplvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gjt2z4 <= 1'b1;
  else
    Gjt2z4 <= Iplvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ukt2z4 <= 1'b1;
  else
    Ukt2z4 <= Bplvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Imt2z4 <= 1'b1;
  else
    Imt2z4 <= Uolvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wnt2z4 <= 1'b1;
  else
    Wnt2z4 <= Bilvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lpt2z4 <= 1'b1;
  else
    Lpt2z4 <= Fdlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Art2z4 <= 1'b1;
  else
    Art2z4 <= Q8lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pst2z4 <= 1'b1;
  else
    Pst2z4 <= B4lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eut2z4 <= 1'b1;
  else
    Eut2z4 <= Mzkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tvt2z4 <= 1'b1;
  else
    Tvt2z4 <= Evkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ixt2z4 <= 1'b1;
  else
    Ixt2z4 <= Pqkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wyt2z4 <= 1'b1;
  else
    Wyt2z4 <= Amkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K0u2z4 <= 1'b1;
  else
    K0u2z4 <= Lhkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y1u2z4 <= 1'b1;
  else
    Y1u2z4 <= Wckvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M3u2z4 <= 1'b1;
  else
    M3u2z4 <= A8kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B5u2z4 <= 1'b1;
  else
    B5u2z4 <= L3kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q6u2z4 <= 1'b1;
  else
    Q6u2z4 <= Hujvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F8u2z4 <= 1'b1;
  else
    F8u2z4 <= Spjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U9u2z4 <= 1'b1;
  else
    U9u2z4 <= Dljvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jbu2z4 <= 1'b1;
  else
    Jbu2z4 <= Ogjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ycu2z4 <= 1'b1;
  else
    Ycu2z4 <= Zbjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Neu2z4 <= 1'b1;
  else
    Neu2z4 <= K7jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cgu2z4 <= 1'b1;
  else
    Cgu2z4 <= V2jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rhu2z4 <= 1'b1;
  else
    Rhu2z4 <= Rtivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gju2z4 <= 1'b1;
  else
    Gju2z4 <= Cpivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uku2z4 <= 1'b1;
  else
    Uku2z4 <= Nkivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Imu2z4 <= 1'b1;
  else
    Imu2z4 <= Yfivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wnu2z4 <= 1'b1;
  else
    Wnu2z4 <= Jbivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lpu2z4 <= 1'b1;
  else
    Lpu2z4 <= Enlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aru2z4 <= 1'b1;
  else
    Aru2z4 <= Xmlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Psu2z4 <= 1'b1;
  else
    Psu2z4 <= Qmlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Duu2z4 <= 1'b1;
  else
    Duu2z4 <= Jmlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rvu2z4 <= 1'b1;
  else
    Rvu2z4 <= Cmlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fxu2z4 <= 1'b1;
  else
    Fxu2z4 <= Nhlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uyu2z4 <= 1'b1;
  else
    Uyu2z4 <= Rclvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J0v2z4 <= 1'b1;
  else
    J0v2z4 <= C8lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y1v2z4 <= 1'b1;
  else
    Y1v2z4 <= N3lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N3v2z4 <= 1'b1;
  else
    N3v2z4 <= Yykvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C5v2z4 <= 1'b1;
  else
    C5v2z4 <= Qukvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R6v2z4 <= 1'b1;
  else
    R6v2z4 <= Bqkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F8v2z4 <= 1'b1;
  else
    F8v2z4 <= Mlkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T9v2z4 <= 1'b1;
  else
    T9v2z4 <= Xgkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hbv2z4 <= 1'b1;
  else
    Hbv2z4 <= Ickvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vcv2z4 <= 1'b1;
  else
    Vcv2z4 <= M7kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kev2z4 <= 1'b1;
  else
    Kev2z4 <= X2kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zfv2z4 <= 1'b1;
  else
    Zfv2z4 <= Ttjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ohv2z4 <= 1'b1;
  else
    Ohv2z4 <= Epjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Djv2z4 <= 1'b1;
  else
    Djv2z4 <= Pkjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Skv2z4 <= 1'b1;
  else
    Skv2z4 <= Agjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hmv2z4 <= 1'b1;
  else
    Hmv2z4 <= Lbjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wnv2z4 <= 1'b1;
  else
    Wnv2z4 <= W6jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lpv2z4 <= 1'b1;
  else
    Lpv2z4 <= H2jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Arv2z4 <= 1'b1;
  else
    Arv2z4 <= Dtivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Psv2z4 <= 1'b1;
  else
    Psv2z4 <= Ooivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Duv2z4 <= 1'b1;
  else
    Duv2z4 <= Zjivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rvv2z4 <= 1'b1;
  else
    Rvv2z4 <= Kfivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fxv2z4 <= 1'b1;
  else
    Fxv2z4 <= Vaivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uyv2z4 <= 1'b0;
  else
    Uyv2z4 <= H6mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G0w2z4 <= 1'b1;
  else
    G0w2z4 <= Acnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R1w2z4 <= 1'b1;
  else
    R1w2z4 <= Ocnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C3w2z4 <= 1'b0;
  else
    C3w2z4 <= Ufnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S4w2z4 <= 1'b0;
  else
    S4w2z4 <= Srhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I6w2z4 <= 1'b0;
  else
    I6w2z4 <= X7mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U7w2z4 <= 1'b0;
  else
    U7w2z4 <= Q7mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G9w2z4 <= 1'b1;
  else
    G9w2z4 <= Lrhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vaw2z4 <= 1'b0;
  else
    Vaw2z4 <= Erhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jcw2z4 <= 1'b1;
  else
    Jcw2z4 <= Xqhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ydw2z4 <= 1'b1;
  else
    Ydw2z4 <= Qqhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mfw2z4 <= 1'b1;
  else
    Mfw2z4 <= Jqhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ahw2z4 <= 1'b1;
  else
    Ahw2z4 <= Cqhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Oiw2z4 <= 1'b1;
  else
    Oiw2z4 <= Vphvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ckw2z4 <= 1'b1;
  else
    Ckw2z4 <= Ophvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qlw2z4 <= 1'b1;
  else
    Qlw2z4 <= Hphvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Enw2z4 <= 1'b1;
  else
    Enw2z4 <= Aphvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sow2z4 <= 1'b1;
  else
    Sow2z4 <= Tohvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gqw2z4 <= 1'b1;
  else
    Gqw2z4 <= Mohvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Urw2z4 <= 1'b1;
  else
    Urw2z4 <= Fohvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Itw2z4 <= 1'b1;
  else
    Itw2z4 <= Ynhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xuw2z4 <= 1'b1;
  else
    Xuw2z4 <= Rnhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mww2z4 <= 1'b1;
  else
    Mww2z4 <= Knhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Byw2z4 <= 1'b1;
  else
    Byw2z4 <= Dnhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qzw2z4 <= 1'b1;
  else
    Qzw2z4 <= Wmhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F1x2z4 <= 1'b1;
  else
    F1x2z4 <= Pmhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U2x2z4 <= 1'b1;
  else
    U2x2z4 <= Hjnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J4x2z4 <= 1'b1;
  else
    J4x2z4 <= Imhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U5x2z4 <= 1'b0;
  else
    U5x2z4 <= F5mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G7x2z4 <= 1'b1;
  else
    G7x2z4 <= Bmhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R8x2z4 <= 1'b1;
  else
    R8x2z4 <= Ulhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cax2z4 <= 1'b1;
  else
    Cax2z4 <= Nlhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nbx2z4 <= 1'b1;
  else
    Nbx2z4 <= Glhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ycx2z4 <= 1'b1;
  else
    Ycx2z4 <= Zkhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jex2z4 <= 1'b1;
  else
    Jex2z4 <= Skhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ufx2z4 <= 1'b1;
  else
    Ufx2z4 <= Lkhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fhx2z4 <= 1'b1;
  else
    Fhx2z4 <= Ekhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rix2z4 <= 1'b1;
  else
    Rix2z4 <= Xjhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dkx2z4 <= 1'b1;
  else
    Dkx2z4 <= Qjhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Plx2z4 <= 1'b1;
  else
    Plx2z4 <= Jjhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bnx2z4 <= 1'b1;
  else
    Bnx2z4 <= Cjhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nox2z4 <= 1'b1;
  else
    Nox2z4 <= Vihvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zpx2z4 <= 1'b1;
  else
    Zpx2z4 <= Oihvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lrx2z4 <= 1'b1;
  else
    Lrx2z4 <= Hihvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xsx2z4 <= 1'b1;
  else
    Xsx2z4 <= Aihvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jux2z4 <= 1'b1;
  else
    Jux2z4 <= Thhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vvx2z4 <= 1'b1;
  else
    Vvx2z4 <= Mhhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hxx2z4 <= 1'b1;
  else
    Hxx2z4 <= Fhhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tyx2z4 <= 1'b1;
  else
    Tyx2z4 <= Yghvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F0y2z4 <= 1'b1;
  else
    F0y2z4 <= Yanvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T1y2z4 <= 1'b1;
  else
    T1y2z4 <= Slnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I3y2z4 <= 1'b1;
  else
    I3y2z4 <= Ranvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W4y2z4 <= 1'b1;
  else
    W4y2z4 <= Kanvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K6y2z4 <= 1'b1;
  else
    K6y2z4 <= Danvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y7y2z4 <= 1'b1;
  else
    Y7y2z4 <= W9nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M9y2z4 <= 1'b1;
  else
    M9y2z4 <= P9nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bby2z4 <= 1'b1;
  else
    Bby2z4 <= I9nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qcy2z4 <= 1'b1;
  else
    Qcy2z4 <= B9nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fey2z4 <= 1'b1;
  else
    Fey2z4 <= N8nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ufy2z4 <= 1'b1;
  else
    Ufy2z4 <= G8nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jhy2z4 <= 1'b0;
  else
    Jhy2z4 <= Z7nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Viy2z4 <= 1'b1;
  else
    Viy2z4 <= L7nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jky2z4 <= 1'b1;
  else
    Jky2z4 <= E7nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xly2z4 <= 1'b1;
  else
    Xly2z4 <= X6nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lny2z4 <= 1'b1;
  else
    Lny2z4 <= Q6nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zoy2z4 <= 1'b1;
  else
    Zoy2z4 <= J6nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nqy2z4 <= 1'b1;
  else
    Nqy2z4 <= C6nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bsy2z4 <= 1'b1;
  else
    Bsy2z4 <= V5nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pty2z4 <= 1'b1;
  else
    Pty2z4 <= O5nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dvy2z4 <= 1'b1;
  else
    Dvy2z4 <= H5nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Swy2z4 <= 1'b1;
  else
    Swy2z4 <= A5nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hyy2z4 <= 1'b1;
  else
    Hyy2z4 <= T4nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wzy2z4 <= 1'b1;
  else
    Wzy2z4 <= Rghvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K1z2z4 <= 1'b1;
  else
    K1z2z4 <= I3mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C3z2z4 <= 1'b1;
  else
    C3z2z4 <= B3mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U4z2z4 <= 1'b1;
  else
    U4z2z4 <= Vllvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I6z2z4 <= 1'b1;
  else
    I6z2z4 <= Kghvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W7z2z4 <= 1'b1;
  else
    W7z2z4 <= Dghvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K9z2z4 <= 1'b1;
  else
    K9z2z4 <= Wfhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yaz2z4 <= 1'b1;
  else
    Yaz2z4 <= Pfhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mcz2z4 <= 1'b1;
  else
    Mcz2z4 <= Allvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aez2z4 <= 1'b1;
  else
    Aez2z4 <= Tklvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pfz2z4 <= 1'b1;
  else
    Pfz2z4 <= Mklvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ehz2z4 <= 1'b1;
  else
    Ehz2z4 <= Oslvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tiz2z4 <= 1'b1;
  else
    Tiz2z4 <= Hslvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ikz2z4 <= 1'b1;
  else
    Ikz2z4 <= Aslvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wlz2z4 <= 1'b1;
  else
    Wlz2z4 <= Trlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Knz2z4 <= 1'b1;
  else
    Knz2z4 <= Mrlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yoz2z4 <= 1'b1;
  else
    Yoz2z4 <= Tdlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nqz2z4 <= 1'b1;
  else
    Nqz2z4 <= P4lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Csz2z4 <= 1'b1;
  else
    Csz2z4 <= A0lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rtz2z4 <= 1'b1;
  else
    Rtz2z4 <= Drkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fvz2z4 <= 1'b1;
  else
    Fvz2z4 <= Omkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Twz2z4 <= 1'b1;
  else
    Twz2z4 <= Zhkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hyz2z4 <= 1'b1;
  else
    Hyz2z4 <= Kdkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vzz2z4 <= 1'b1;
  else
    Vzz2z4 <= O8kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K103z4 <= 1'b1;
  else
    K103z4 <= Gqjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z203z4 <= 1'b1;
  else
    Z203z4 <= Rljvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O403z4 <= 1'b1;
  else
    O403z4 <= Chjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D603z4 <= 1'b1;
  else
    D603z4 <= Ncjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S703z4 <= 1'b1;
  else
    S703z4 <= J3jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H903z4 <= 1'b1;
  else
    H903z4 <= Fuivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wa03z4 <= 1'b1;
  else
    Wa03z4 <= Qpivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kc03z4 <= 1'b1;
  else
    Kc03z4 <= Mgivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yd03z4 <= 1'b1;
  else
    Yd03z4 <= Xtlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nf03z4 <= 1'b1;
  else
    Nf03z4 <= Qtlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ch03z4 <= 1'b1;
  else
    Ch03z4 <= Jtlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qi03z4 <= 1'b1;
  else
    Qi03z4 <= Ctlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ek03z4 <= 1'b1;
  else
    Ek03z4 <= Vslvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sl03z4 <= 1'b1;
  else
    Sl03z4 <= Aelvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hn03z4 <= 1'b1;
  else
    Hn03z4 <= W4lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wo03z4 <= 1'b1;
  else
    Wo03z4 <= H0lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lq03z4 <= 1'b1;
  else
    Lq03z4 <= Krkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zr03z4 <= 1'b1;
  else
    Zr03z4 <= Vmkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nt03z4 <= 1'b1;
  else
    Nt03z4 <= Gikvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bv03z4 <= 1'b1;
  else
    Bv03z4 <= Rdkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pw03z4 <= 1'b1;
  else
    Pw03z4 <= V8kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ey03z4 <= 1'b1;
  else
    Ey03z4 <= Nqjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tz03z4 <= 1'b1;
  else
    Tz03z4 <= Yljvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I113z4 <= 1'b1;
  else
    I113z4 <= Jhjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X213z4 <= 1'b1;
  else
    X213z4 <= Ucjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M413z4 <= 1'b1;
  else
    M413z4 <= Q3jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B613z4 <= 1'b1;
  else
    B613z4 <= Muivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q713z4 <= 1'b1;
  else
    Q713z4 <= Xpivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E913z4 <= 1'b1;
  else
    E913z4 <= Tgivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sa13z4 <= 1'b1;
  else
    Sa13z4 <= Gvlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hc13z4 <= 1'b1;
  else
    Hc13z4 <= Zulvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wd13z4 <= 1'b1;
  else
    Wd13z4 <= Sulvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kf13z4 <= 1'b1;
  else
    Kf13z4 <= Lulvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yg13z4 <= 1'b1;
  else
    Yg13z4 <= Eulvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mi13z4 <= 1'b1;
  else
    Mi13z4 <= Ghlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bk13z4 <= 1'b1;
  else
    Bk13z4 <= Kclvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ql13z4 <= 1'b1;
  else
    Ql13z4 <= V7lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fn13z4 <= 1'b1;
  else
    Fn13z4 <= G3lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uo13z4 <= 1'b1;
  else
    Uo13z4 <= Rykvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jq13z4 <= 1'b1;
  else
    Jq13z4 <= Jukvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yr13z4 <= 1'b1;
  else
    Yr13z4 <= Upkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mt13z4 <= 1'b1;
  else
    Mt13z4 <= Flkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Av13z4 <= 1'b1;
  else
    Av13z4 <= Qgkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ow13z4 <= 1'b1;
  else
    Ow13z4 <= Bckvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cy13z4 <= 1'b1;
  else
    Cy13z4 <= F7kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rz13z4 <= 1'b1;
  else
    Rz13z4 <= Q2kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G123z4 <= 1'b1;
  else
    G123z4 <= Mtjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V223z4 <= 1'b1;
  else
    V223z4 <= Xojvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K423z4 <= 1'b1;
  else
    K423z4 <= Ikjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z523z4 <= 1'b1;
  else
    Z523z4 <= Tfjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O723z4 <= 1'b1;
  else
    O723z4 <= Ebjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D923z4 <= 1'b1;
  else
    D923z4 <= P6jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sa23z4 <= 1'b1;
  else
    Sa23z4 <= A2jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hc23z4 <= 1'b1;
  else
    Hc23z4 <= Wsivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wd23z4 <= 1'b1;
  else
    Wd23z4 <= Hoivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kf23z4 <= 1'b1;
  else
    Kf23z4 <= Sjivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yg23z4 <= 1'b1;
  else
    Yg23z4 <= Dfivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mi23z4 <= 1'b1;
  else
    Mi23z4 <= Oaivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bk23z4 <= 1'b1;
  else
    Bk23z4 <= Pwlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ql23z4 <= 1'b1;
  else
    Ql23z4 <= Iwlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fn23z4 <= 1'b1;
  else
    Fn23z4 <= Bwlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    To23z4 <= 1'b1;
  else
    To23z4 <= Uvlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hq23z4 <= 1'b1;
  else
    Hq23z4 <= Nvlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vr23z4 <= 1'b1;
  else
    Vr23z4 <= Zglvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kt23z4 <= 1'b1;
  else
    Kt23z4 <= Dclvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zu23z4 <= 1'b1;
  else
    Zu23z4 <= O7lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ow23z4 <= 1'b1;
  else
    Ow23z4 <= Z2lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dy23z4 <= 1'b1;
  else
    Dy23z4 <= Kykvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sz23z4 <= 1'b1;
  else
    Sz23z4 <= Cukvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H133z4 <= 1'b1;
  else
    H133z4 <= Npkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V233z4 <= 1'b1;
  else
    V233z4 <= Ykkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J433z4 <= 1'b1;
  else
    J433z4 <= Jgkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X533z4 <= 1'b1;
  else
    X533z4 <= Ubkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L733z4 <= 1'b1;
  else
    L733z4 <= Y6kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A933z4 <= 1'b1;
  else
    A933z4 <= J2kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pa33z4 <= 1'b1;
  else
    Pa33z4 <= Ftjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ec33z4 <= 1'b1;
  else
    Ec33z4 <= Qojvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Td33z4 <= 1'b1;
  else
    Td33z4 <= Bkjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    If33z4 <= 1'b1;
  else
    If33z4 <= Mfjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xg33z4 <= 1'b1;
  else
    Xg33z4 <= Xajvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mi33z4 <= 1'b1;
  else
    Mi33z4 <= I6jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bk33z4 <= 1'b1;
  else
    Bk33z4 <= T1jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ql33z4 <= 1'b1;
  else
    Ql33z4 <= Psivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fn33z4 <= 1'b1;
  else
    Fn33z4 <= Aoivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    To33z4 <= 1'b1;
  else
    To33z4 <= Ljivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hq33z4 <= 1'b1;
  else
    Hq33z4 <= Weivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vr33z4 <= 1'b1;
  else
    Vr33z4 <= Haivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kt33z4 <= 1'b1;
  else
    Kt33z4 <= Yxlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zu33z4 <= 1'b1;
  else
    Zu33z4 <= Rxlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ow33z4 <= 1'b1;
  else
    Ow33z4 <= Kxlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cy33z4 <= 1'b1;
  else
    Cy33z4 <= Dxlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qz33z4 <= 1'b1;
  else
    Qz33z4 <= Wwlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E143z4 <= 1'b1;
  else
    E143z4 <= Sglvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T243z4 <= 1'b1;
  else
    T243z4 <= Wblvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I443z4 <= 1'b1;
  else
    I443z4 <= H7lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X543z4 <= 1'b1;
  else
    X543z4 <= S2lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M743z4 <= 1'b1;
  else
    M743z4 <= Dykvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B943z4 <= 1'b1;
  else
    B943z4 <= Vtkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qa43z4 <= 1'b1;
  else
    Qa43z4 <= Gpkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ec43z4 <= 1'b1;
  else
    Ec43z4 <= Rkkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sd43z4 <= 1'b1;
  else
    Sd43z4 <= Cgkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gf43z4 <= 1'b1;
  else
    Gf43z4 <= Nbkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ug43z4 <= 1'b1;
  else
    Ug43z4 <= R6kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ji43z4 <= 1'b1;
  else
    Ji43z4 <= C2kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yj43z4 <= 1'b1;
  else
    Yj43z4 <= Ysjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nl43z4 <= 1'b1;
  else
    Nl43z4 <= Jojvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cn43z4 <= 1'b1;
  else
    Cn43z4 <= Ujjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ro43z4 <= 1'b1;
  else
    Ro43z4 <= Ffjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gq43z4 <= 1'b1;
  else
    Gq43z4 <= Qajvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vr43z4 <= 1'b1;
  else
    Vr43z4 <= B6jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kt43z4 <= 1'b1;
  else
    Kt43z4 <= M1jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zu43z4 <= 1'b1;
  else
    Zu43z4 <= Isivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ow43z4 <= 1'b1;
  else
    Ow43z4 <= Tnivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cy43z4 <= 1'b1;
  else
    Cy43z4 <= Ejivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qz43z4 <= 1'b1;
  else
    Qz43z4 <= Peivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E153z4 <= 1'b1;
  else
    E153z4 <= Aaivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T253z4 <= 1'b1;
  else
    T253z4 <= Hzlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I453z4 <= 1'b1;
  else
    I453z4 <= Azlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X553z4 <= 1'b1;
  else
    X553z4 <= Tylvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L753z4 <= 1'b1;
  else
    L753z4 <= Mylvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z853z4 <= 1'b1;
  else
    Z853z4 <= Fylvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Na53z4 <= 1'b1;
  else
    Na53z4 <= Lglvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cc53z4 <= 1'b1;
  else
    Cc53z4 <= Pblvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rd53z4 <= 1'b1;
  else
    Rd53z4 <= A7lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gf53z4 <= 1'b1;
  else
    Gf53z4 <= L2lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vg53z4 <= 1'b1;
  else
    Vg53z4 <= Wxkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ki53z4 <= 1'b1;
  else
    Ki53z4 <= Otkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zj53z4 <= 1'b1;
  else
    Zj53z4 <= Zokvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nl53z4 <= 1'b1;
  else
    Nl53z4 <= Kkkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bn53z4 <= 1'b1;
  else
    Bn53z4 <= Vfkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Po53z4 <= 1'b1;
  else
    Po53z4 <= Gbkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dq53z4 <= 1'b1;
  else
    Dq53z4 <= K6kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sr53z4 <= 1'b1;
  else
    Sr53z4 <= V1kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ht53z4 <= 1'b1;
  else
    Ht53z4 <= Rsjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wu53z4 <= 1'b1;
  else
    Wu53z4 <= Cojvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lw53z4 <= 1'b1;
  else
    Lw53z4 <= Njjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ay53z4 <= 1'b1;
  else
    Ay53z4 <= Yejvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pz53z4 <= 1'b1;
  else
    Pz53z4 <= Jajvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E163z4 <= 1'b1;
  else
    E163z4 <= U5jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T263z4 <= 1'b1;
  else
    T263z4 <= F1jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I463z4 <= 1'b1;
  else
    I463z4 <= Bsivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X563z4 <= 1'b1;
  else
    X563z4 <= Mnivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L763z4 <= 1'b1;
  else
    L763z4 <= Xiivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z863z4 <= 1'b1;
  else
    Z863z4 <= Ieivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Na63z4 <= 1'b1;
  else
    Na63z4 <= T9ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cc63z4 <= 1'b1;
  else
    Cc63z4 <= Q0mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rd63z4 <= 1'b1;
  else
    Rd63z4 <= J0mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gf63z4 <= 1'b1;
  else
    Gf63z4 <= C0mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ug63z4 <= 1'b1;
  else
    Ug63z4 <= Vzlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ii63z4 <= 1'b1;
  else
    Ii63z4 <= Ozlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wj63z4 <= 1'b1;
  else
    Wj63z4 <= Eglvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ll63z4 <= 1'b1;
  else
    Ll63z4 <= Iblvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    An63z4 <= 1'b1;
  else
    An63z4 <= T6lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Po63z4 <= 1'b1;
  else
    Po63z4 <= E2lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eq63z4 <= 1'b1;
  else
    Eq63z4 <= Pxkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tr63z4 <= 1'b1;
  else
    Tr63z4 <= Htkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    It63z4 <= 1'b1;
  else
    It63z4 <= Sokvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wu63z4 <= 1'b1;
  else
    Wu63z4 <= Dkkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kw63z4 <= 1'b1;
  else
    Kw63z4 <= Ofkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yx63z4 <= 1'b1;
  else
    Yx63z4 <= Zakvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mz63z4 <= 1'b1;
  else
    Mz63z4 <= D6kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B173z4 <= 1'b1;
  else
    B173z4 <= O1kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q273z4 <= 1'b1;
  else
    Q273z4 <= Ksjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F473z4 <= 1'b1;
  else
    F473z4 <= Vnjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U573z4 <= 1'b1;
  else
    U573z4 <= Gjjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J773z4 <= 1'b1;
  else
    J773z4 <= Rejvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y873z4 <= 1'b1;
  else
    Y873z4 <= Cajvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Na73z4 <= 1'b1;
  else
    Na73z4 <= N5jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cc73z4 <= 1'b1;
  else
    Cc73z4 <= Y0jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rd73z4 <= 1'b1;
  else
    Rd73z4 <= Urivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gf73z4 <= 1'b1;
  else
    Gf73z4 <= Fnivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ug73z4 <= 1'b1;
  else
    Ug73z4 <= Qiivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ii73z4 <= 1'b1;
  else
    Ii73z4 <= Beivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wj73z4 <= 1'b1;
  else
    Wj73z4 <= M9ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ll73z4 <= 1'b1;
  else
    Ll73z4 <= Z1mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    An73z4 <= 1'b1;
  else
    An73z4 <= S1mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Po73z4 <= 1'b1;
  else
    Po73z4 <= L1mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dq73z4 <= 1'b1;
  else
    Dq73z4 <= E1mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rr73z4 <= 1'b1;
  else
    Rr73z4 <= X0mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ft73z4 <= 1'b1;
  else
    Ft73z4 <= Xflvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uu73z4 <= 1'b1;
  else
    Uu73z4 <= Bblvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jw73z4 <= 1'b1;
  else
    Jw73z4 <= M6lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yx73z4 <= 1'b1;
  else
    Yx73z4 <= X1lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nz73z4 <= 1'b1;
  else
    Nz73z4 <= Ixkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C183z4 <= 1'b1;
  else
    C183z4 <= Atkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R283z4 <= 1'b1;
  else
    R283z4 <= Lokvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F483z4 <= 1'b1;
  else
    F483z4 <= Wjkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T583z4 <= 1'b1;
  else
    T583z4 <= Hfkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H783z4 <= 1'b1;
  else
    H783z4 <= Sakvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V883z4 <= 1'b1;
  else
    V883z4 <= W5kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ka83z4 <= 1'b1;
  else
    Ka83z4 <= H1kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zb83z4 <= 1'b1;
  else
    Zb83z4 <= Dsjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Od83z4 <= 1'b1;
  else
    Od83z4 <= Onjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Df83z4 <= 1'b1;
  else
    Df83z4 <= Zijvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sg83z4 <= 1'b1;
  else
    Sg83z4 <= Kejvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hi83z4 <= 1'b1;
  else
    Hi83z4 <= V9jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wj83z4 <= 1'b1;
  else
    Wj83z4 <= G5jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ll83z4 <= 1'b1;
  else
    Ll83z4 <= R0jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    An83z4 <= 1'b1;
  else
    An83z4 <= Nrivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Po83z4 <= 1'b1;
  else
    Po83z4 <= Ymivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dq83z4 <= 1'b1;
  else
    Dq83z4 <= Jiivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rr83z4 <= 1'b1;
  else
    Rr83z4 <= Udivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ft83z4 <= 1'b1;
  else
    Ft83z4 <= F9ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uu83z4 <= 1'b1;
  else
    Uu83z4 <= Jflvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jw83z4 <= 1'b1;
  else
    Jw83z4 <= Nalvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yx83z4 <= 1'b1;
  else
    Yx83z4 <= Y5lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nz83z4 <= 1'b1;
  else
    Nz83z4 <= J1lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C193z4 <= 1'b1;
  else
    C193z4 <= Uwkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    R293z4 <= 1'b1;
  else
    R293z4 <= Mskvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G493z4 <= 1'b1;
  else
    G493z4 <= Xnkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U593z4 <= 1'b1;
  else
    U593z4 <= Fskvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I793z4 <= 1'b1;
  else
    I793z4 <= Pgnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W893z4 <= 1'b1;
  else
    W893z4 <= Ijkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ka93z4 <= 1'b1;
  else
    Ka93z4 <= Tekvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yb93z4 <= 1'b1;
  else
    Yb93z4 <= Eakvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Md93z4 <= 1'b1;
  else
    Md93z4 <= I5kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bf93z4 <= 1'b1;
  else
    Bf93z4 <= T0kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qg93z4 <= 1'b1;
  else
    Qg93z4 <= Prjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fi93z4 <= 1'b1;
  else
    Fi93z4 <= Anjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uj93z4 <= 1'b1;
  else
    Uj93z4 <= Lijvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jl93z4 <= 1'b1;
  else
    Jl93z4 <= Wdjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ym93z4 <= 1'b1;
  else
    Ym93z4 <= Eijvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    No93z4 <= 1'b1;
  else
    No93z4 <= H9jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cq93z4 <= 1'b1;
  else
    Cq93z4 <= S4jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rr93z4 <= 1'b1;
  else
    Rr93z4 <= D0jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gt93z4 <= 1'b1;
  else
    Gt93z4 <= Zqivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vu93z4 <= 1'b1;
  else
    Vu93z4 <= Kmivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jw93z4 <= 1'b1;
  else
    Jw93z4 <= K4mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xx93z4 <= 1'b1;
  else
    Xx93z4 <= Mekvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lz93z4 <= 1'b0;
  else
    Lz93z4 <= Jknvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B1a3z4 <= 1'b0;
  else
    B1a3z4 <= Hdmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P2a3z4 <= 1'b0;
  else
    P2a3z4 <= Admvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D4a3z4 <= 1'b1;
  else
    D4a3z4 <= Ivmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U5a3z4 <= 1'b1;
  else
    U5a3z4 <= Pvmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    L7a3z4 <= 1'b1;
  else
    L7a3z4 <= Dwmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C9a3z4 <= 1'b1;
  else
    C9a3z4 <= Rwmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Taa3z4 <= 1'b1;
  else
    Taa3z4 <= Hymvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jca3z4 <= 1'b1;
  else
    Jca3z4 <= Umnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aea3z4 <= 1'b1;
  else
    Aea3z4 <= Jzmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qfa3z4 <= 1'b1;
  else
    Qfa3z4 <= Czmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gha3z4 <= 1'b1;
  else
    Gha3z4 <= Vymvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wia3z4 <= 1'b1;
  else
    Wia3z4 <= Oymvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mka3z4 <= 1'b1;
  else
    Mka3z4 <= Aymvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cma3z4 <= 1'b1;
  else
    Cma3z4 <= Ltmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tna3z4 <= 1'b0;
  else
    Tna3z4 <= Xzmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jpa3z4 <= 1'b1;
  else
    Jpa3z4 <= Bomvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ara3z4 <= 1'b1;
  else
    Ara3z4 <= Dpmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rsa3z4 <= 1'b1;
  else
    Rsa3z4 <= Kpmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Iua3z4 <= 1'b1;
  else
    Iua3z4 <= Ypmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zva3z4 <= 1'b1;
  else
    Zva3z4 <= Mqmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qxa3z4 <= 1'b1;
  else
    Qxa3z4 <= Vrmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gza3z4 <= 1'b1;
  else
    Gza3z4 <= Csmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W0b3z4 <= 1'b1;
  else
    W0b3z4 <= Jsmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M2b3z4 <= 1'b1;
  else
    M2b3z4 <= Qsmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C4b3z4 <= 1'b1;
  else
    C4b3z4 <= Xsmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S5b3z4 <= 1'b0;
  else
    S5b3z4 <= Qzmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J7b3z4 <= 1'b1;
  else
    J7b3z4 <= Txmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z8b3z4 <= 1'b1;
  else
    Z8b3z4 <= Ormvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pab3z4 <= 1'b0;
  else
    Pab3z4 <= Smmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gcb3z4 <= 1'b0;
  else
    Gcb3z4 <= Okmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xdb3z4 <= 1'b0;
  else
    Xdb3z4 <= Kimvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nfb3z4 <= 1'b1;
  else
    Nfb3z4 <= Mxmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dhb3z4 <= 1'b1;
  else
    Dhb3z4 <= Hrmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tib3z4 <= 1'b0;
  else
    Tib3z4 <= Lmmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kkb3z4 <= 1'b0;
  else
    Kkb3z4 <= Hkmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bmb3z4 <= 1'b0;
  else
    Bmb3z4 <= Dimvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rnb3z4 <= 1'b0;
  else
    Rnb3z4 <= S8mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ipb3z4 <= 1'b0;
  else
    Ipb3z4 <= R1ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zqb3z4 <= 1'b0;
  else
    Zqb3z4 <= Gmnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qsb3z4 <= 1'b0;
  else
    Qsb3z4 <= Iamvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hub3z4 <= 1'b0;
  else
    Hub3z4 <= Y1ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Yvb3z4 <= 1'b0;
  else
    Yvb3z4 <= Bamvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pxb3z4 <= 1'b0;
  else
    Pxb3z4 <= F2ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gzb3z4 <= 1'b0;
  else
    Gzb3z4 <= N9mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X0c3z4 <= 1'b0;
  else
    X0c3z4 <= W0ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O2c3z4 <= 1'b0;
  else
    O2c3z4 <= G9mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F4c3z4 <= 1'b0;
  else
    F4c3z4 <= D1ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W5c3z4 <= 1'b0;
  else
    W5c3z4 <= Z8mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N7c3z4 <= 1'b0;
  else
    N7c3z4 <= K1ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E9c3z4 <= 1'b0;
  else
    E9c3z4 <= Y4mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vac3z4 <= 1'b0;
  else
    Vac3z4 <= M2ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mcc3z4 <= 1'b0;
  else
    Mcc3z4 <= E0nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bec3z4 <= 1'b0;
  else
    Bec3z4 <= L0nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qfc3z4 <= 1'b0;
  else
    Qfc3z4 <= S0nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fhc3z4 <= 1'b0;
  else
    Fhc3z4 <= Z0nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uic3z4 <= 1'b0;
  else
    Uic3z4 <= G1nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jkc3z4 <= 1'b0;
  else
    Jkc3z4 <= N1nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ylc3z4 <= 1'b0;
  else
    Ylc3z4 <= U1nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nnc3z4 <= 1'b0;
  else
    Nnc3z4 <= P2nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dpc3z4 <= 1'b0;
  else
    Dpc3z4 <= D3nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tqc3z4 <= 1'b0;
  else
    Tqc3z4 <= R3nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jsc3z4 <= 1'b0;
  else
    Jsc3z4 <= Y3nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ztc3z4 <= 1'b0;
  else
    Ztc3z4 <= Cknvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ovc3z4 <= 1'b1;
  else
    Ovc3z4 <= Bjkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cxc3z4 <= 1'b1;
  else
    Cxc3z4 <= Vhivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qyc3z4 <= 1'b1;
  else
    Qyc3z4 <= Gdivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    E0d3z4 <= 1'b1;
  else
    E0d3z4 <= R8ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T1d3z4 <= 1'b1;
  else
    T1d3z4 <= Ifhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H3d3z4 <= 1'b1;
  else
    H3d3z4 <= G2mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    V4d3z4 <= 1'b1;
  else
    V4d3z4 <= Bfhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    G6d3z4 <= 1'b1;
  else
    G6d3z4 <= Sqivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T7d3z4 <= 1'b0;
  else
    T7d3z4 <= Lfmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J9d3z4 <= 1'b0;
  else
    J9d3z4 <= Ggmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zad3z4 <= 1'b0;
  else
    Zad3z4 <= Zfmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pcd3z4 <= 1'b0;
  else
    Pcd3z4 <= Sfmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fed3z4 <= 1'b0;
  else
    Fed3z4 <= Efmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vfd3z4 <= 1'b0;
  else
    Vfd3z4 <= Xemvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lhd3z4 <= 1'b0;
  else
    Lhd3z4 <= Qemvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bjd3z4 <= 1'b0;
  else
    Bjd3z4 <= Jemvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rkd3z4 <= 1'b1;
  else
    Rkd3z4 <= Hvivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gmd3z4 <= 1'b1;
  else
    Gmd3z4 <= Uehvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Snd3z4 <= 1'b1;
  else
    Snd3z4 <= Ovivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hpd3z4 <= 1'b1;
  else
    Hpd3z4 <= Vvivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wqd3z4 <= 1'b1;
  else
    Wqd3z4 <= Cwivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lsd3z4 <= 1'b1;
  else
    Lsd3z4 <= Jwivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aud3z4 <= 1'b1;
  else
    Aud3z4 <= Qwivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pvd3z4 <= 1'b1;
  else
    Pvd3z4 <= Xwivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Exd3z4 <= 1'b1;
  else
    Exd3z4 <= Exivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tyd3z4 <= 1'b1;
  else
    Tyd3z4 <= Lxivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I0e3z4 <= 1'b1;
  else
    I0e3z4 <= Sxivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    X1e3z4 <= 1'b1;
  else
    X1e3z4 <= Zxivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M3e3z4 <= 1'b1;
  else
    M3e3z4 <= Gyivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B5e3z4 <= 1'b1;
  else
    B5e3z4 <= Nyivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q6e3z4 <= 1'b1;
  else
    Q6e3z4 <= Uyivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    F8e3z4 <= 1'b1;
  else
    F8e3z4 <= Bzivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    U9e3z4 <= 1'b1;
  else
    U9e3z4 <= Izivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ibe3z4 <= 1'b1;
  else
    Ibe3z4 <= Pzivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wce3z4 <= 1'b1;
  else
    Wce3z4 <= Wzivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lee3z4 <= 1'b0;
  else
    Lee3z4 <= W2nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bge3z4 <= 1'b1;
  else
    Bge3z4 <= Kwmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    She3z4 <= 1'b1;
  else
    She3z4 <= Fqmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jje3z4 <= 1'b0;
  else
    Jje3z4 <= J7mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ble3z4 <= 1'b0;
  else
    Ble3z4 <= Uzhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tme3z4 <= 1'b1;
  else
    Tme3z4 <= Nehvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Foe3z4 <= 1'b1;
  else
    Foe3z4 <= Gehvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rpe3z4 <= 1'b1;
  else
    Rpe3z4 <= Blivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fre3z4 <= 1'b1;
  else
    Fre3z4 <= Ilivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tse3z4 <= 1'b1;
  else
    Tse3z4 <= Plivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hue3z4 <= 1'b1;
  else
    Hue3z4 <= Wlivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vve3z4 <= 1'b0;
  else
    Vve3z4 <= I2nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kxe3z4 <= 1'b1;
  else
    Kxe3z4 <= Ywmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aze3z4 <= 1'b1;
  else
    Aze3z4 <= Tqmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q0f3z4 <= 1'b0;
  else
    Q0f3z4 <= V6mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    H2f3z4 <= 1'b0;
  else
    H2f3z4 <= B2nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    W3f3z4 <= 1'b1;
  else
    W3f3z4 <= Fxmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M5f3z4 <= 1'b1;
  else
    M5f3z4 <= Armvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    C7f3z4 <= 1'b0;
  else
    C7f3z4 <= O6mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T8f3z4 <= 1'b0;
  else
    T8f3z4 <= P0ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kaf3z4 <= 1'b1;
  else
    Kaf3z4 <= Zdhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wbf3z4 <= 1'b1;
  else
    Wbf3z4 <= C4ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ldf3z4 <= 1'b1;
  else
    Ldf3z4 <= Q4ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aff3z4 <= 1'b1;
  else
    Aff3z4 <= X4ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pgf3z4 <= 1'b1;
  else
    Pgf3z4 <= E5ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eif3z4 <= 1'b1;
  else
    Eif3z4 <= L5ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tjf3z4 <= 1'b1;
  else
    Tjf3z4 <= S5ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ilf3z4 <= 1'b1;
  else
    Ilf3z4 <= Z5ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xmf3z4 <= 1'b1;
  else
    Xmf3z4 <= G6ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Mof3z4 <= 1'b1;
  else
    Mof3z4 <= N6ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Bqf3z4 <= 1'b1;
  else
    Bqf3z4 <= U6ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qrf3z4 <= 1'b1;
  else
    Qrf3z4 <= I7ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ftf3z4 <= 1'b1;
  else
    Ftf3z4 <= P7ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uuf3z4 <= 1'b1;
  else
    Uuf3z4 <= D8ivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Jwf3z4 <= 1'b1;
  else
    Jwf3z4 <= Sdhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vxf3z4 <= 1'b1;
  else
    Vxf3z4 <= Y7jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kzf3z4 <= 1'b1;
  else
    Kzf3z4 <= F8jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z0g3z4 <= 1'b1;
  else
    Z0g3z4 <= M8jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    O2g3z4 <= 1'b1;
  else
    O2g3z4 <= T8jvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    D4g3z4 <= 1'b0;
  else
    D4g3z4 <= K3nvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    T5g3z4 <= 1'b1;
  else
    T5g3z4 <= Wvmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    K7g3z4 <= 1'b1;
  else
    K7g3z4 <= Rpmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B9g3z4 <= 1'b1;
  else
    B9g3z4 <= Ldhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Nag3z4 <= 1'b1;
  else
    Nag3z4 <= Ewjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ccg3z4 <= 1'b1;
  else
    Ccg3z4 <= Lwjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rdg3z4 <= 1'b1;
  else
    Rdg3z4 <= Swjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Gfg3z4 <= 1'b1;
  else
    Gfg3z4 <= Zwjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Vgg3z4 <= 1'b1;
  else
    Vgg3z4 <= Gxjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Kig3z4 <= 1'b1;
  else
    Kig3z4 <= Nxjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zjg3z4 <= 1'b1;
  else
    Zjg3z4 <= Uxjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Olg3z4 <= 1'b1;
  else
    Olg3z4 <= Byjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Dng3z4 <= 1'b1;
  else
    Dng3z4 <= Iyjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Sog3z4 <= 1'b1;
  else
    Sog3z4 <= Pyjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hqg3z4 <= 1'b1;
  else
    Hqg3z4 <= Wyjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wrg3z4 <= 1'b1;
  else
    Wrg3z4 <= Dzjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ltg3z4 <= 1'b1;
  else
    Ltg3z4 <= Kzjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Avg3z4 <= 1'b1;
  else
    Avg3z4 <= Rzjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Pwg3z4 <= 1'b1;
  else
    Pwg3z4 <= Yzjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Eyg3z4 <= 1'b1;
  else
    Eyg3z4 <= F0kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tzg3z4 <= 1'b1;
  else
    Tzg3z4 <= M0kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I1h3z4 <= 1'b1;
  else
    I1h3z4 <= Ztmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Z2h3z4 <= 1'b1;
  else
    Z2h3z4 <= Unmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Q4h3z4 <= 1'b0;
  else
    Q4h3z4 <= R4mvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    I6h3z4 <= 1'b0;
  else
    I6h3z4 <= Kbmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    A8h3z4 <= 1'b1;
  else
    A8h3z4 <= Z3kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    P9h3z4 <= 1'b1;
  else
    P9h3z4 <= G4kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ebh3z4 <= 1'b1;
  else
    Ebh3z4 <= N4kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tch3z4 <= 1'b1;
  else
    Tch3z4 <= U4kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ieh3z4 <= 1'b1;
  else
    Ieh3z4 <= Stmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Zfh3z4 <= 1'b1;
  else
    Zfh3z4 <= Q9kvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ohh3z4 <= 1'b1;
  else
    Ohh3z4 <= Khnvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Djh3z4 <= 1'b1;
  else
    Djh3z4 <= E9lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Skh3z4 <= 1'b1;
  else
    Skh3z4 <= L9lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Hmh3z4 <= 1'b1;
  else
    Hmh3z4 <= S9lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Wnh3z4 <= 1'b1;
  else
    Wnh3z4 <= Z9lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lph3z4 <= 1'b1;
  else
    Lph3z4 <= Xbivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Arh3z4 <= 1'b1;
  else
    Arh3z4 <= Ecivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Psh3z4 <= 1'b1;
  else
    Psh3z4 <= Lcivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Euh3z4 <= 1'b1;
  else
    Euh3z4 <= Scivx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Tvh3z4 <= 1'b1;
  else
    Tvh3z4 <= Vujvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ixh3z4 <= 1'b1;
  else
    Ixh3z4 <= Cvjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Xyh3z4 <= 1'b1;
  else
    Xyh3z4 <= Jvjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    M0i3z4 <= 1'b1;
  else
    M0i3z4 <= Qvjvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    B2i3z4 <= 1'b1;
  else
    B2i3z4 <= Uumvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    S3i3z4 <= 1'b1;
  else
    S3i3z4 <= Pomvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    J5i3z4 <= 1'b1;
  else
    J5i3z4 <= Pilvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Y6i3z4 <= 1'b1;
  else
    Y6i3z4 <= Wilvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    N8i3z4 <= 1'b1;
  else
    N8i3z4 <= Djlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Cai3z4 <= 1'b1;
  else
    Cai3z4 <= Kjlvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Rbi3z4 <= 1'b1;
  else
    Rbi3z4 <= Edhvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ddi3z4 <= 1'b1;
  else
    Ddi3z4 <= Gnmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Uei3z4 <= 1'b1;
  else
    Uei3z4 <= Zmmvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Lgi3z4 <= 1'b1;
  else
    Lgi3z4 <= C1lvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Aii3z4 <= 1'b0;
  else
    Aii3z4 <= Xchvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Qji3z4 <= 1'b1;
  else
    Qji3z4 <= Svkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Fli3z4 <= 1'b1;
  else
    Fli3z4 <= Zvkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Umi3z4 <= 1'b1;
  else
    Umi3z4 <= Gwkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Joi3z4 <= 1'b1;
  else
    Joi3z4 <= Nwkvx4;

always @(posedge hclk or negedge hreset_n)
  if(~hreset_n)
    Ypi3z4 <= 1'b0;
  else
    Ypi3z4 <= Qchvx4;

endmodule

//------------------------------------------------------------------------------
// EOF
//------------------------------------------------------------------------------

